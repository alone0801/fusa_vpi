
//__CDS_SVN_TAG__
// $URL: file:///projects/cdnsfs/svn_repo/ifss_vmgr_flow_proj/trunk/demo/SRC/NL/dut.mapped.no_escapes.v $ $Id: dut.mapped.no_escapes.v 667 2016-11-15 17:44:59Z ferlini $
// ------------------------------------------------------------------------------
// Copyright (c) 2016 by Cadence Design Systems, All Rights Reserved.
//
// This software is provided as is without warranty of any kind.  The entire risk
// as to the results and performance of this software is assumed by the user.
//
// Cadence Design Systems disclaims all warranties, either express or implied,
// including but not limited, the implied warranties of merchantability, fitness
// for a particular purpose, title and no infringement, with respect to this
// software.
//
// No technical support is guaranteed for this code. If you have any suggestion
// or improvement feel free to contact your Cadence representative.
// ------------------------------------------------------------------------------
//__CDS_SVN_TAG__

// Generated by Cadence Encounter(R) RTL Compiler RC14.23 - v14.20-s027_1

// Verification Directory fv/dut 

module crc_gen_DATA_WIDTH32_POLYNOMIAL_BITS8(clk, rst_n, data_in,
     crc_val);
  input clk, rst_n;
  input [31:0] data_in;
  output [7:0] crc_val;
  wire clk, rst_n;
  wire [31:0] data_in;
  wire [7:0] crc_val;
  wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7;
  wire n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15;
  wire n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23;
  wire n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31;
  wire n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39;
  wire n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47;
  wire n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55;
  wire n_56, n_57, n_58, n_60, n_61, n_67, n_68;
  XNOR2X1 g1048(.A (n_30), .B (n_67), .Y (crc_val[0]));
  XOR2XL g1049(.A (n_48), .B (n_68), .Y (crc_val[3]));
  XNOR2X1 g1050(.A (data_in[10]), .B (n_60), .Y (n_68));
  XNOR2X1 g1051(.A (data_in[22]), .B (n_60), .Y (n_67));
  CLKXOR2X1 g1052(.A (n_29), .B (n_61), .Y (crc_val[4]));
  XNOR2X1 g1053(.A (n_52), .B (n_58), .Y (crc_val[7]));
  XNOR2X1 g1054(.A (n_39), .B (n_51), .Y (crc_val[5]));
  XNOR2X1 g1055(.A (n_38), .B (n_54), .Y (crc_val[1]));
  CLKXOR2X1 g1056(.A (n_28), .B (n_53), .Y (crc_val[6]));
  XNOR2X1 g1057(.A (n_21), .B (n_55), .Y (n_61));
  XNOR2X1 g1058(.A (n_42), .B (n_57), .Y (n_60));
  CLKXOR2X1 g1059(.A (n_40), .B (n_56), .Y (crc_val[2]));
  XNOR2X1 g1060(.A (n_30), .B (n_49), .Y (n_58));
  XNOR2X1 g1061(.A (n_13), .B (n_47), .Y (n_57));
  XNOR2X1 g1062(.A (n_3), .B (n_46), .Y (n_56));
  XNOR2X1 g1063(.A (data_in[10]), .B (n_50), .Y (n_55));
  XNOR2X1 g1064(.A (data_in[21]), .B (n_50), .Y (n_54));
  XNOR2X1 g1065(.A (n_19), .B (n_45), .Y (n_53));
  XNOR2X1 g1066(.A (n_20), .B (n_44), .Y (n_52));
  XNOR2X1 g1067(.A (n_34), .B (n_49), .Y (n_51));
  XNOR2X1 g1068(.A (n_27), .B (n_43), .Y (n_50));
  XNOR2X1 g1069(.A (data_in[11]), .B (n_36), .Y (n_49));
  XNOR2X1 g1070(.A (n_16), .B (n_41), .Y (n_48));
  XNOR2X1 g1071(.A (data_in[0]), .B (n_36), .Y (n_47));
  XNOR2X1 g1072(.A (data_in[24]), .B (n_37), .Y (n_46));
  XNOR2X1 g1073(.A (n_10), .B (n_37), .Y (n_45));
  XNOR2X1 g1074(.A (data_in[30]), .B (n_41), .Y (n_44));
  XNOR2X1 g1075(.A (n_18), .B (n_32), .Y (n_43));
  XNOR2X1 g1076(.A (n_12), .B (n_35), .Y (n_42));
  XNOR2X1 g1077(.A (n_1), .B (n_33), .Y (n_41));
  XNOR2X1 g1078(.A (n_11), .B (n_34), .Y (n_40));
  XNOR2X1 g1079(.A (n_9), .B (n_31), .Y (n_39));
  XNOR2X1 g1080(.A (n_22), .B (n_35), .Y (n_38));
  XNOR2X1 g1081(.A (n_17), .B (n_26), .Y (n_37));
  XNOR2X1 g1082(.A (n_14), .B (n_25), .Y (n_36));
  XNOR2X1 g1083(.A (data_in[17]), .B (n_10), .Y (n_33));
  XNOR2X1 g1084(.A (data_in[30]), .B (n_11), .Y (n_32));
  XNOR2X1 g1085(.A (data_in[24]), .B (n_2), .Y (n_35));
  XNOR2X1 g1086(.A (data_in[18]), .B (n_8), .Y (n_31));
  XNOR2X1 g1087(.A (data_in[17]), .B (n_0), .Y (n_34));
  XNOR2X1 g1088(.A (n_7), .B (n_12), .Y (n_29));
  XNOR2X1 g1089(.A (n_5), .B (n_24), .Y (n_30));
  XNOR2X1 g1090(.A (n_23), .B (n_24), .Y (n_28));
  XNOR2X1 g1091(.A (n_6), .B (n_8), .Y (n_27));
  XNOR2X1 g1092(.A (n_15), .B (n_9), .Y (n_26));
  XNOR2X1 g1093(.A (n_4), .B (n_23), .Y (n_25));
  XNOR2X1 g1094(.A (data_in[23]), .B (data_in[18]), .Y (n_22));
  XNOR2X1 g1095(.A (data_in[2]), .B (data_in[18]), .Y (n_24));
  XNOR2X1 g1096(.A (data_in[27]), .B (data_in[17]), .Y (n_21));
  XNOR2X1 g1097(.A (data_in[24]), .B (data_in[0]), .Y (n_20));
  XNOR2X1 g1098(.A (data_in[29]), .B (data_in[10]), .Y (n_19));
  XNOR2X1 g1099(.A (data_in[16]), .B (data_in[0]), .Y (n_18));
  XNOR2X1 g1100(.A (data_in[19]), .B (data_in[16]), .Y (n_17));
  XNOR2X1 g1101(.A (data_in[16]), .B (data_in[9]), .Y (n_16));
  XNOR2X1 g1102(.A (data_in[22]), .B (data_in[21]), .Y (n_15));
  XNOR2X1 g1103(.A (data_in[31]), .B (data_in[21]), .Y (n_14));
  XNOR2X1 g1104(.A (data_in[28]), .B (data_in[12]), .Y (n_23));
  XNOR2X1 g1105(.A (data_in[29]), .B (data_in[13]), .Y (n_13));
  XNOR2X1 g1106(.A (data_in[3]), .B (data_in[19]), .Y (n_12));
  XNOR2X1 g1107(.A (data_in[26]), .B (data_in[11]), .Y (n_7));
  XNOR2X1 g1108(.A (data_in[12]), .B (data_in[14]), .Y (n_6));
  XNOR2X1 g1109(.A (data_in[26]), .B (data_in[25]), .Y (n_5));
  XNOR2X1 g1110(.A (data_in[8]), .B (data_in[31]), .Y (n_11));
  XNOR2X1 g1111(.A (data_in[27]), .B (data_in[1]), .Y (n_4));
  XNOR2X1 g1112(.A (data_in[6]), .B (data_in[14]), .Y (n_10));
  XNOR2X1 g1113(.A (data_in[5]), .B (data_in[13]), .Y (n_9));
  XNOR2X1 g1114(.A (data_in[1]), .B (data_in[25]), .Y (n_3));
  XNOR2X1 g1115(.A (data_in[7]), .B (data_in[15]), .Y (n_2));
  XNOR2X1 g1116(.A (data_in[23]), .B (data_in[20]), .Y (n_1));
  XNOR2X1 g1117(.A (data_in[4]), .B (data_in[20]), .Y (n_8));
  XNOR2X1 g1118(.A (data_in[15]), .B (data_in[9]), .Y (n_0));
endmodule

module crc_chk_DATA_WIDTH32_POLYNOMIAL_BITS8(clk, rst_n, data_in,
     crc_in, data_out, err_detected, err_corrected);
  input clk, rst_n;
  input [31:0] data_in;
  input [7:0] crc_in;
  output [31:0] data_out;
  output err_detected, err_corrected;
  wire clk, rst_n;
  wire [31:0] data_in;
  wire [7:0] crc_in;
  wire [31:0] data_out;
  wire err_detected, err_corrected;
  wire [7:0] crc_calc;
  wire UNCONNECTED_HIER_Z, UNCONNECTED_HIER_Z0, n_0, n_1, n_2, n_3,
       n_4, n_5;
  wire n_6, n_7, n_8, n_9, n_10, n_11, n_12, n_13;
  wire n_14, n_15, n_16, n_17;
  crc_gen_DATA_WIDTH32_POLYNOMIAL_BITS8 crc_gen_i(.clk
       (UNCONNECTED_HIER_Z), .rst_n (UNCONNECTED_HIER_Z0), .data_in
       (data_in), .crc_val (crc_calc));
  DFFRHQX1 err_detected_reg(.RN (rst_n), .CK (clk), .D (n_17), .Q
       (err_detected));
  NAND2X1 g318(.A (n_10), .B (n_16), .Y (n_17));
  AOI221X1 g319(.A0 (crc_in[4]), .A1 (n_2), .B0 (crc_in[6]), .B1 (n_1),
       .C0 (n_15), .Y (n_16));
  OAI211X1 g320(.A0 (crc_in[6]), .A1 (n_1), .B0 (n_9), .C0 (n_14), .Y
       (n_15));
  NOR4X1 g321(.A (n_8), .B (n_7), .C (n_12), .D (n_13), .Y (n_14));
  OAI221X1 g322(.A0 (crc_in[3]), .A1 (n_4), .B0 (crc_in[4]), .B1 (n_2),
       .C0 (n_11), .Y (n_13));
  OAI222X1 g323(.A0 (n_3), .A1 (crc_calc[2]), .B0 (crc_in[0]), .B1
       (n_5), .C0 (crc_in[2]), .C1 (n_0), .Y (n_12));
  AOI22X1 g324(.A0 (crc_in[3]), .A1 (n_4), .B0 (n_6), .B1
       (crc_calc[1]), .Y (n_11));
  XNOR2X1 g325(.A (crc_in[7]), .B (crc_calc[7]), .Y (n_10));
  XNOR2X1 g326(.A (crc_in[5]), .B (crc_calc[5]), .Y (n_9));
  NOR2X1 g327(.A (n_6), .B (crc_calc[1]), .Y (n_8));
  NOR2BX1 g328(.AN (crc_in[0]), .B (crc_calc[0]), .Y (n_7));
  INVX1 g329(.A (crc_in[1]), .Y (n_6));
  INVX1 g330(.A (crc_calc[0]), .Y (n_5));
  INVX1 g331(.A (crc_calc[3]), .Y (n_4));
  INVX1 g332(.A (crc_in[2]), .Y (n_3));
  INVX1 g333(.A (crc_calc[4]), .Y (n_2));
  INVX1 g334(.A (crc_calc[6]), .Y (n_1));
  INVX1 g335(.A (crc_calc[2]), .Y (n_0));
endmodule

module crc_gen_DATA_WIDTH32_POLYNOMIAL_BITS8_2(clk, rst_n, data_in,
     crc_val);
  input clk, rst_n;
  input [31:0] data_in;
  output [7:0] crc_val;
  wire clk, rst_n;
  wire [31:0] data_in;
  wire [7:0] crc_val;
  wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7;
  wire n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15;
  wire n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23;
  wire n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31;
  wire n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39;
  wire n_40, n_41, n_42, n_43, n_44, n_45, n_46, n_47;
  wire n_48, n_49, n_50, n_51, n_52, n_53, n_54, n_55;
  wire n_56, n_57, n_58, n_59, n_61, n_62, n_68, n_69;
  XNOR2X1 g1081(.A (n_30), .B (n_68), .Y (crc_val[0]));
  XOR2XL g1082(.A (n_49), .B (n_69), .Y (crc_val[3]));
  XNOR2X1 g1083(.A (data_in[10]), .B (n_61), .Y (n_69));
  XNOR2X1 g1084(.A (data_in[22]), .B (n_61), .Y (n_68));
  XOR2XL g1085(.A (n_31), .B (n_62), .Y (crc_val[4]));
  XNOR2X1 g1086(.A (n_52), .B (n_58), .Y (crc_val[7]));
  XNOR2X1 g1087(.A (n_44), .B (n_59), .Y (crc_val[5]));
  XNOR2X1 g1088(.A (n_39), .B (n_54), .Y (crc_val[1]));
  XOR2XL g1089(.A (n_28), .B (n_53), .Y (crc_val[6]));
  XNOR2X1 g1090(.A (n_22), .B (n_55), .Y (n_62));
  XNOR2X1 g1091(.A (n_41), .B (n_57), .Y (n_61));
  XOR2XL g1092(.A (n_40), .B (n_56), .Y (crc_val[2]));
  XNOR2X1 g1093(.A (n_11), .B (n_50), .Y (n_59));
  XNOR2X1 g1094(.A (n_30), .B (n_50), .Y (n_58));
  XNOR2X1 g1095(.A (n_15), .B (n_48), .Y (n_57));
  XNOR2X1 g1096(.A (n_6), .B (n_47), .Y (n_56));
  XNOR2X1 g1097(.A (data_in[10]), .B (n_51), .Y (n_55));
  XNOR2X1 g1098(.A (data_in[21]), .B (n_51), .Y (n_54));
  XNOR2X1 g1099(.A (n_20), .B (n_46), .Y (n_53));
  XNOR2X1 g1100(.A (n_21), .B (n_45), .Y (n_52));
  XNOR2X1 g1101(.A (n_27), .B (n_43), .Y (n_51));
  XNOR2X1 g1102(.A (data_in[11]), .B (n_36), .Y (n_50));
  XNOR2X1 g1103(.A (n_17), .B (n_42), .Y (n_49));
  XNOR2X1 g1104(.A (data_in[0]), .B (n_36), .Y (n_48));
  XNOR2X1 g1105(.A (data_in[24]), .B (n_37), .Y (n_47));
  XNOR2X1 g1106(.A (n_8), .B (n_37), .Y (n_46));
  XNOR2X1 g1107(.A (data_in[30]), .B (n_42), .Y (n_45));
  XNOR2X1 g1108(.A (n_14), .B (n_38), .Y (n_44));
  XNOR2X1 g1109(.A (n_19), .B (n_34), .Y (n_43));
  XNOR2X1 g1110(.A (n_3), .B (n_35), .Y (n_42));
  XNOR2X1 g1111(.A (n_10), .B (n_33), .Y (n_41));
  XNOR2X1 g1112(.A (n_9), .B (n_32), .Y (n_40));
  XNOR2X1 g1113(.A (n_23), .B (n_33), .Y (n_39));
  XNOR2X1 g1114(.A (data_in[13]), .B (n_32), .Y (n_38));
  XNOR2X1 g1115(.A (n_18), .B (n_26), .Y (n_37));
  XNOR2X1 g1116(.A (n_24), .B (n_29), .Y (n_36));
  XNOR2X1 g1117(.A (data_in[17]), .B (n_8), .Y (n_35));
  XNOR2X1 g1118(.A (data_in[30]), .B (n_9), .Y (n_34));
  XNOR2X1 g1119(.A (data_in[24]), .B (n_2), .Y (n_33));
  XNOR2X1 g1120(.A (data_in[17]), .B (n_0), .Y (n_32));
  XNOR2X1 g1121(.A (n_7), .B (n_10), .Y (n_31));
  XNOR2X1 g1122(.A (n_4), .B (n_25), .Y (n_30));
  XNOR2X1 g1123(.A (n_1), .B (n_12), .Y (n_29));
  XNOR2X1 g1124(.A (n_12), .B (n_25), .Y (n_28));
  XNOR2X1 g1125(.A (n_5), .B (n_11), .Y (n_27));
  XNOR2X1 g1126(.A (n_16), .B (n_13), .Y (n_26));
  XNOR2X1 g1127(.A (data_in[2]), .B (data_in[18]), .Y (n_25));
  XNOR2X1 g1128(.A (data_in[21]), .B (data_in[31]), .Y (n_24));
  XNOR2X1 g1129(.A (data_in[18]), .B (data_in[23]), .Y (n_23));
  XNOR2X1 g1130(.A (data_in[17]), .B (data_in[27]), .Y (n_22));
  XNOR2X1 g1131(.A (data_in[0]), .B (data_in[24]), .Y (n_21));
  XNOR2X1 g1132(.A (data_in[10]), .B (data_in[29]), .Y (n_20));
  XNOR2X1 g1133(.A (data_in[0]), .B (data_in[16]), .Y (n_19));
  XNOR2X1 g1134(.A (data_in[16]), .B (data_in[19]), .Y (n_18));
  XNOR2X1 g1135(.A (data_in[9]), .B (data_in[16]), .Y (n_17));
  XNOR2X1 g1136(.A (data_in[21]), .B (data_in[22]), .Y (n_16));
  XNOR2X1 g1137(.A (data_in[13]), .B (data_in[29]), .Y (n_15));
  XNOR2X1 g1138(.A (data_in[5]), .B (data_in[18]), .Y (n_14));
  XNOR2X1 g1139(.A (data_in[5]), .B (data_in[13]), .Y (n_13));
  XNOR2X1 g1140(.A (data_in[12]), .B (data_in[28]), .Y (n_12));
  XNOR2X1 g1141(.A (data_in[4]), .B (data_in[20]), .Y (n_11));
  XNOR2X1 g1142(.A (data_in[3]), .B (data_in[19]), .Y (n_10));
  XNOR2X1 g1143(.A (data_in[11]), .B (data_in[26]), .Y (n_7));
  XNOR2X1 g1144(.A (data_in[1]), .B (data_in[25]), .Y (n_6));
  XNOR2X1 g1145(.A (data_in[12]), .B (data_in[14]), .Y (n_5));
  XNOR2X1 g1146(.A (data_in[25]), .B (data_in[26]), .Y (n_4));
  XNOR2X1 g1147(.A (data_in[8]), .B (data_in[31]), .Y (n_9));
  XNOR2X1 g1148(.A (data_in[6]), .B (data_in[14]), .Y (n_8));
  XNOR2X1 g1149(.A (data_in[20]), .B (data_in[23]), .Y (n_3));
  XNOR2X1 g1150(.A (data_in[7]), .B (data_in[15]), .Y (n_2));
  XNOR2X1 g1151(.A (data_in[1]), .B (data_in[27]), .Y (n_1));
  XNOR2X1 g1152(.A (data_in[9]), .B (data_in[15]), .Y (n_0));
endmodule

module mem_with_crc_DATA_WIDTH32_POLYNOMIAL_BITS8(clk, rst_n, mem_wr,
     mem_data_in, crc_data_in, mem_data_out, crc_data_out);
  input clk, rst_n, mem_wr;
  input [31:0] mem_data_in;
  input [7:0] crc_data_in;
  output [31:0] mem_data_out;
  output [7:0] crc_data_out;
  wire clk, rst_n, mem_wr;
  wire [31:0] mem_data_in;
  wire [7:0] crc_data_in;
  wire [31:0] mem_data_out;
  wire [7:0] crc_data_out;
  wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7;
  wire n_8, n_9, n_10, n_11, n_12, n_13, n_14, n_15;
  wire n_16, n_17, n_18, n_19, n_20, n_21, n_22, n_23;
  wire n_24, n_25, n_26, n_27, n_28, n_29, n_30, n_31;
  wire n_32, n_33, n_34, n_35, n_36, n_37, n_38, n_39;
  DFFRHQX1 mem_crc_reg_0(.RN (rst_n), .CK (clk), .D (n_31), .Q
       (crc_data_out[0]));
  DFFRHQX1 mem_crc_reg_1(.RN (rst_n), .CK (clk), .D (n_24), .Q
       (crc_data_out[1]));
  DFFRHQX1 mem_reg_10(.RN (rst_n), .CK (clk), .D (n_0), .Q
       (mem_data_out[10]));
  DFFRHQX1 mem_reg_11(.RN (rst_n), .CK (clk), .D (n_39), .Q
       (mem_data_out[11]));
  DFFRHQX1 mem_reg_12(.RN (rst_n), .CK (clk), .D (n_38), .Q
       (mem_data_out[12]));
  DFFRHQX1 mem_reg_13(.RN (rst_n), .CK (clk), .D (n_37), .Q
       (mem_data_out[13]));
  DFFRHQX1 mem_reg_14(.RN (rst_n), .CK (clk), .D (n_36), .Q
       (mem_data_out[14]));
  DFFRHQX1 mem_reg_15(.RN (rst_n), .CK (clk), .D (n_35), .Q
       (mem_data_out[15]));
  DFFRHQX1 mem_reg_16(.RN (rst_n), .CK (clk), .D (n_34), .Q
       (mem_data_out[16]));
  DFFRHQX1 mem_reg_17(.RN (rst_n), .CK (clk), .D (n_33), .Q
       (mem_data_out[17]));
  DFFRHQX1 mem_reg_18(.RN (rst_n), .CK (clk), .D (n_32), .Q
       (mem_data_out[18]));
  DFFRHQX1 mem_reg_19(.RN (rst_n), .CK (clk), .D (n_30), .Q
       (mem_data_out[19]));
  DFFRHQX1 mem_reg_2(.RN (rst_n), .CK (clk), .D (n_29), .Q
       (mem_data_out[2]));
  DFFRHQX1 mem_reg_20(.RN (rst_n), .CK (clk), .D (n_28), .Q
       (mem_data_out[20]));
  DFFRHQX1 mem_reg_21(.RN (rst_n), .CK (clk), .D (n_27), .Q
       (mem_data_out[21]));
  DFFRHQX1 mem_reg_22(.RN (rst_n), .CK (clk), .D (n_25), .Q
       (mem_data_out[22]));
  DFFRHQX1 mem_reg_23(.RN (rst_n), .CK (clk), .D (n_23), .Q
       (mem_data_out[23]));
  DFFRHQX1 mem_reg_24(.RN (rst_n), .CK (clk), .D (n_21), .Q
       (mem_data_out[24]));
  DFFRHQX1 mem_crc_reg_2(.RN (rst_n), .CK (clk), .D (n_22), .Q
       (crc_data_out[2]));
  DFFRHQX1 mem_crc_reg_3(.RN (rst_n), .CK (clk), .D (n_18), .Q
       (crc_data_out[3]));
  DFFRHQX1 mem_reg_25(.RN (rst_n), .CK (clk), .D (n_20), .Q
       (mem_data_out[25]));
  DFFRHQX1 mem_reg_26(.RN (rst_n), .CK (clk), .D (n_19), .Q
       (mem_data_out[26]));
  DFFRHQX1 mem_reg_27(.RN (rst_n), .CK (clk), .D (n_17), .Q
       (mem_data_out[27]));
  DFFRHQX1 mem_reg_28(.RN (rst_n), .CK (clk), .D (n_15), .Q
       (mem_data_out[28]));
  DFFRHQX1 mem_crc_reg_4(.RN (rst_n), .CK (clk), .D (n_16), .Q
       (crc_data_out[4]));
  DFFRHQX1 mem_reg_29(.RN (rst_n), .CK (clk), .D (n_14), .Q
       (mem_data_out[29]));
  DFFRHQX1 mem_reg_3(.RN (rst_n), .CK (clk), .D (n_12), .Q
       (mem_data_out[3]));
  DFFRHQX1 mem_crc_reg_5(.RN (rst_n), .CK (clk), .D (n_13), .Q
       (crc_data_out[5]));
  DFFRHQX1 mem_reg_30(.RN (rst_n), .CK (clk), .D (n_11), .Q
       (mem_data_out[30]));
  DFFRHQX1 mem_reg_31(.RN (rst_n), .CK (clk), .D (n_9), .Q
       (mem_data_out[31]));
  DFFRHQX1 mem_crc_reg_6(.RN (rst_n), .CK (clk), .D (n_10), .Q
       (crc_data_out[6]));
  DFFRHQX1 mem_crc_reg_7(.RN (rst_n), .CK (clk), .D (n_5), .Q
       (crc_data_out[7]));
  DFFRHQX1 mem_reg_4(.RN (rst_n), .CK (clk), .D (n_8), .Q
       (mem_data_out[4]));
  DFFRHQX1 mem_reg_5(.RN (rst_n), .CK (clk), .D (n_7), .Q
       (mem_data_out[5]));
  DFFRHQX1 mem_reg_6(.RN (rst_n), .CK (clk), .D (n_6), .Q
       (mem_data_out[6]));
  DFFRHQX1 mem_reg_7(.RN (rst_n), .CK (clk), .D (n_26), .Q
       (mem_data_out[7]));
  DFFRHQX1 mem_reg_0(.RN (rst_n), .CK (clk), .D (n_4), .Q
       (mem_data_out[0]));
  DFFRHQX1 mem_reg_8(.RN (rst_n), .CK (clk), .D (n_3), .Q
       (mem_data_out[8]));
  DFFRHQX1 mem_reg_9(.RN (rst_n), .CK (clk), .D (n_1), .Q
       (mem_data_out[9]));
  DFFRHQX1 mem_reg_1(.RN (rst_n), .CK (clk), .D (n_2), .Q
       (mem_data_out[1]));
  MX2XL g84(.A (mem_data_out[11]), .B (mem_data_in[11]), .S0 (mem_wr),
       .Y (n_39));
  MX2XL g85(.A (mem_data_out[12]), .B (mem_data_in[12]), .S0 (mem_wr),
       .Y (n_38));
  MX2XL g86(.A (mem_data_out[13]), .B (mem_data_in[13]), .S0 (mem_wr),
       .Y (n_37));
  MX2XL g87(.A (mem_data_out[14]), .B (mem_data_in[14]), .S0 (mem_wr),
       .Y (n_36));
  MX2XL g88(.A (mem_data_out[15]), .B (mem_data_in[15]), .S0 (mem_wr),
       .Y (n_35));
  MX2XL g89(.A (mem_data_out[16]), .B (mem_data_in[16]), .S0 (mem_wr),
       .Y (n_34));
  MX2XL g90(.A (mem_data_out[17]), .B (mem_data_in[17]), .S0 (mem_wr),
       .Y (n_33));
  MX2XL g91(.A (mem_data_out[18]), .B (mem_data_in[18]), .S0 (mem_wr),
       .Y (n_32));
  MX2XL g92(.A (crc_data_out[0]), .B (crc_data_in[0]), .S0 (mem_wr), .Y
       (n_31));
  MX2XL g93(.A (mem_data_out[19]), .B (mem_data_in[19]), .S0 (mem_wr),
       .Y (n_30));
  MX2XL g94(.A (mem_data_out[2]), .B (mem_data_in[2]), .S0 (mem_wr), .Y
       (n_29));
  MX2XL g95(.A (mem_data_out[20]), .B (mem_data_in[20]), .S0 (mem_wr),
       .Y (n_28));
  MX2XL g96(.A (mem_data_out[21]), .B (mem_data_in[21]), .S0 (mem_wr),
       .Y (n_27));
  MX2XL g97(.A (mem_data_out[7]), .B (mem_data_in[7]), .S0 (mem_wr), .Y
       (n_26));
  MX2XL g98(.A (mem_data_out[22]), .B (mem_data_in[22]), .S0 (mem_wr),
       .Y (n_25));
  MX2XL g99(.A (crc_data_out[1]), .B (crc_data_in[1]), .S0 (mem_wr), .Y
       (n_24));
  MX2XL g100(.A (mem_data_out[23]), .B (mem_data_in[23]), .S0 (mem_wr),
       .Y (n_23));
  MX2XL g101(.A (crc_data_out[2]), .B (crc_data_in[2]), .S0 (mem_wr),
       .Y (n_22));
  MX2XL g102(.A (mem_data_out[24]), .B (mem_data_in[24]), .S0 (mem_wr),
       .Y (n_21));
  MX2XL g103(.A (mem_data_out[25]), .B (mem_data_in[25]), .S0 (mem_wr),
       .Y (n_20));
  MX2XL g104(.A (mem_data_out[26]), .B (mem_data_in[26]), .S0 (mem_wr),
       .Y (n_19));
  MX2XL g105(.A (crc_data_out[3]), .B (crc_data_in[3]), .S0 (mem_wr),
       .Y (n_18));
  MX2XL g106(.A (mem_data_out[27]), .B (mem_data_in[27]), .S0 (mem_wr),
       .Y (n_17));
  MX2XL g107(.A (crc_data_out[4]), .B (crc_data_in[4]), .S0 (mem_wr),
       .Y (n_16));
  MX2XL g108(.A (mem_data_out[28]), .B (mem_data_in[28]), .S0 (mem_wr),
       .Y (n_15));
  MX2XL g109(.A (mem_data_out[29]), .B (mem_data_in[29]), .S0 (mem_wr),
       .Y (n_14));
  MX2XL g110(.A (crc_data_out[5]), .B (crc_data_in[5]), .S0 (mem_wr),
       .Y (n_13));
  MX2XL g111(.A (mem_data_out[3]), .B (mem_data_in[3]), .S0 (mem_wr),
       .Y (n_12));
  MX2XL g112(.A (mem_data_out[30]), .B (mem_data_in[30]), .S0 (mem_wr),
       .Y (n_11));
  MX2XL g113(.A (crc_data_out[6]), .B (crc_data_in[6]), .S0 (mem_wr),
       .Y (n_10));
  MX2XL g114(.A (mem_data_out[31]), .B (mem_data_in[31]), .S0 (mem_wr),
       .Y (n_9));
  MX2XL g115(.A (mem_data_out[4]), .B (mem_data_in[4]), .S0 (mem_wr),
       .Y (n_8));
  MX2XL g116(.A (mem_data_out[5]), .B (mem_data_in[5]), .S0 (mem_wr),
       .Y (n_7));
  MX2XL g117(.A (mem_data_out[6]), .B (mem_data_in[6]), .S0 (mem_wr),
       .Y (n_6));
  MX2XL g118(.A (crc_data_out[7]), .B (crc_data_in[7]), .S0 (mem_wr),
       .Y (n_5));
  MX2XL g119(.A (mem_data_out[0]), .B (mem_data_in[0]), .S0 (mem_wr),
       .Y (n_4));
  MX2XL g120(.A (mem_data_out[8]), .B (mem_data_in[8]), .S0 (mem_wr),
       .Y (n_3));
  MX2XL g121(.A (mem_data_out[1]), .B (mem_data_in[1]), .S0 (mem_wr),
       .Y (n_2));
  MX2XL g122(.A (mem_data_out[9]), .B (mem_data_in[9]), .S0 (mem_wr),
       .Y (n_1));
  MX2XL g123(.A (mem_data_out[10]), .B (mem_data_in[10]), .S0 (mem_wr),
       .Y (n_0));
endmodule

module crc_mem_DATA_WIDTH32_POLYNOMIAL_BITS8_OUTPUT_FF1(clk, rst_n,
     mem_wr, mem_data_in, mem_data_out, err_detected, err_corrected);
  input clk, rst_n, mem_wr;
  input [31:0] mem_data_in;
  output [31:0] mem_data_out;
  output err_detected, err_corrected;
  wire clk, rst_n, mem_wr;
  wire [31:0] mem_data_in;
  wire [31:0] mem_data_out;
  wire err_detected, err_corrected;
  wire [31:0] mem;
  wire [7:0] mem_crc;
  wire [7:0] crc_wr;
  wire UNCONNECTED, UNCONNECTED0, UNCONNECTED1, UNCONNECTED2,
       UNCONNECTED3, UNCONNECTED4, UNCONNECTED5, UNCONNECTED6;
  wire UNCONNECTED7, UNCONNECTED8, UNCONNECTED9, UNCONNECTED10,
       UNCONNECTED11, UNCONNECTED12, UNCONNECTED13, UNCONNECTED14;
  wire UNCONNECTED15, UNCONNECTED16, UNCONNECTED17, UNCONNECTED18,
       UNCONNECTED19, UNCONNECTED20, UNCONNECTED21, UNCONNECTED22;
  wire UNCONNECTED23, UNCONNECTED24, UNCONNECTED25, UNCONNECTED26,
       UNCONNECTED27, UNCONNECTED28, UNCONNECTED29, UNCONNECTED30;
  wire UNCONNECTED31, UNCONNECTED_HIER_Z1, UNCONNECTED_HIER_Z2;
  crc_chk_DATA_WIDTH32_POLYNOMIAL_BITS8 crc_chk_i(.clk (clk), .rst_n
       (rst_n), .data_in (mem), .crc_in (mem_crc), .data_out
       ({UNCONNECTED30, UNCONNECTED29, UNCONNECTED28, UNCONNECTED27,
       UNCONNECTED26, UNCONNECTED25, UNCONNECTED24, UNCONNECTED23,
       UNCONNECTED22, UNCONNECTED21, UNCONNECTED20, UNCONNECTED19,
       UNCONNECTED18, UNCONNECTED17, UNCONNECTED16, UNCONNECTED15,
       UNCONNECTED14, UNCONNECTED13, UNCONNECTED12, UNCONNECTED11,
       UNCONNECTED10, UNCONNECTED9, UNCONNECTED8, UNCONNECTED7,
       UNCONNECTED6, UNCONNECTED5, UNCONNECTED4, UNCONNECTED3,
       UNCONNECTED2, UNCONNECTED1, UNCONNECTED0, UNCONNECTED}),
       .err_detected (err_detected), .err_corrected (UNCONNECTED31));
  crc_gen_DATA_WIDTH32_POLYNOMIAL_BITS8_2 crc_gen_wr_i(.clk
       (UNCONNECTED_HIER_Z1), .rst_n (UNCONNECTED_HIER_Z2), .data_in
       (mem_data_in), .crc_val (crc_wr));
  mem_with_crc_DATA_WIDTH32_POLYNOMIAL_BITS8 mem_with_crc_i(.clk (clk),
       .rst_n (rst_n), .mem_wr (mem_wr), .mem_data_in (mem_data_in),
       .crc_data_in (crc_wr), .mem_data_out (mem), .crc_data_out
       (mem_crc));
  DFFRHQX1 mem_data_ff_tmp_reg_31(.RN (rst_n), .CK (clk), .D (mem[31]),
       .Q (mem_data_out[31]));
  DFFRHQX1 mem_data_ff_tmp_reg_30(.RN (rst_n), .CK (clk), .D (mem[30]),
       .Q (mem_data_out[30]));
  DFFRHQX1 mem_data_ff_tmp_reg_29(.RN (rst_n), .CK (clk), .D (mem[29]),
       .Q (mem_data_out[29]));
  DFFRHQX1 mem_data_ff_tmp_reg_28(.RN (rst_n), .CK (clk), .D (mem[28]),
       .Q (mem_data_out[28]));
  DFFRHQX1 mem_data_ff_tmp_reg_27(.RN (rst_n), .CK (clk), .D (mem[27]),
       .Q (mem_data_out[27]));
  DFFRHQX1 mem_data_ff_tmp_reg_26(.RN (rst_n), .CK (clk), .D (mem[26]),
       .Q (mem_data_out[26]));
  DFFRHQX1 mem_data_ff_tmp_reg_25(.RN (rst_n), .CK (clk), .D (mem[25]),
       .Q (mem_data_out[25]));
  DFFRHQX1 mem_data_ff_tmp_reg_24(.RN (rst_n), .CK (clk), .D (mem[24]),
       .Q (mem_data_out[24]));
  DFFRHQX1 mem_data_ff_tmp_reg_23(.RN (rst_n), .CK (clk), .D (mem[23]),
       .Q (mem_data_out[23]));
  DFFRHQX1 mem_data_ff_tmp_reg_22(.RN (rst_n), .CK (clk), .D (mem[22]),
       .Q (mem_data_out[22]));
  DFFRHQX1 mem_data_ff_tmp_reg_21(.RN (rst_n), .CK (clk), .D (mem[21]),
       .Q (mem_data_out[21]));
  DFFRHQX1 mem_data_ff_tmp_reg_20(.RN (rst_n), .CK (clk), .D (mem[20]),
       .Q (mem_data_out[20]));
  DFFRHQX1 mem_data_ff_tmp_reg_19(.RN (rst_n), .CK (clk), .D (mem[19]),
       .Q (mem_data_out[19]));
  DFFRHQX1 mem_data_ff_tmp_reg_18(.RN (rst_n), .CK (clk), .D (mem[18]),
       .Q (mem_data_out[18]));
  DFFRHQX1 mem_data_ff_tmp_reg_17(.RN (rst_n), .CK (clk), .D (mem[17]),
       .Q (mem_data_out[17]));
  DFFRHQX1 mem_data_ff_tmp_reg_16(.RN (rst_n), .CK (clk), .D (mem[16]),
       .Q (mem_data_out[16]));
  DFFRHQX1 mem_data_ff_tmp_reg_15(.RN (rst_n), .CK (clk), .D (mem[15]),
       .Q (mem_data_out[15]));
  DFFRHQX1 mem_data_ff_tmp_reg_14(.RN (rst_n), .CK (clk), .D (mem[14]),
       .Q (mem_data_out[14]));
  DFFRHQX1 mem_data_ff_tmp_reg_13(.RN (rst_n), .CK (clk), .D (mem[13]),
       .Q (mem_data_out[13]));
  DFFRHQX1 mem_data_ff_tmp_reg_12(.RN (rst_n), .CK (clk), .D (mem[12]),
       .Q (mem_data_out[12]));
  DFFRHQX1 mem_data_ff_tmp_reg_11(.RN (rst_n), .CK (clk), .D (mem[11]),
       .Q (mem_data_out[11]));
  DFFRHQX1 mem_data_ff_tmp_reg_10(.RN (rst_n), .CK (clk), .D (mem[10]),
       .Q (mem_data_out[10]));
  DFFRHQX1 mem_data_ff_tmp_reg_9(.RN (rst_n), .CK (clk), .D (mem[9]),
       .Q (mem_data_out[9]));
  DFFRHQX1 mem_data_ff_tmp_reg_8(.RN (rst_n), .CK (clk), .D (mem[8]),
       .Q (mem_data_out[8]));
  DFFRHQX1 mem_data_ff_tmp_reg_7(.RN (rst_n), .CK (clk), .D (mem[7]),
       .Q (mem_data_out[7]));
  DFFRHQX1 mem_data_ff_tmp_reg_6(.RN (rst_n), .CK (clk), .D (mem[6]),
       .Q (mem_data_out[6]));
  DFFRHQX1 mem_data_ff_tmp_reg_5(.RN (rst_n), .CK (clk), .D (mem[5]),
       .Q (mem_data_out[5]));
  DFFRHQX1 mem_data_ff_tmp_reg_4(.RN (rst_n), .CK (clk), .D (mem[4]),
       .Q (mem_data_out[4]));
  DFFRHQX1 mem_data_ff_tmp_reg_3(.RN (rst_n), .CK (clk), .D (mem[3]),
       .Q (mem_data_out[3]));
  DFFRHQX1 mem_data_ff_tmp_reg_2(.RN (rst_n), .CK (clk), .D (mem[2]),
       .Q (mem_data_out[2]));
  DFFRHQX1 mem_data_ff_tmp_reg_1(.RN (rst_n), .CK (clk), .D (mem[1]),
       .Q (mem_data_out[1]));
  DFFRHQX1 mem_data_ff_tmp_reg_0(.RN (rst_n), .CK (clk), .D (mem[0]),
       .Q (mem_data_out[0]));
endmodule

module crc_gen_DATA_WIDTH8_POLYNOMIAL_BITS4(clk, rst_n, data_in,
     crc_val);
  input clk, rst_n;
  input [7:0] data_in;
  output [3:0] crc_val;
  wire clk, rst_n;
  wire [7:0] data_in;
  wire [3:0] crc_val;
  wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_8;
  XNOR2X1 g143(.A (n_6), .B (crc_val[0]), .Y (crc_val[1]));
  XNOR2X1 g144(.A (n_5), .B (n_6), .Y (crc_val[2]));
  CLKXOR2X1 g145(.A (data_in[0]), .B (n_8), .Y (crc_val[0]));
  XNOR2X1 g146(.A (n_0), .B (n_4), .Y (n_8));
  CLKXOR2X1 g147(.A (n_4), .B (n_5), .Y (crc_val[3]));
  XNOR2X1 g148(.A (data_in[1]), .B (n_3), .Y (n_6));
  XNOR2X1 g149(.A (data_in[2]), .B (n_2), .Y (n_5));
  XNOR2X1 g150(.A (data_in[3]), .B (n_1), .Y (n_4));
  XNOR2X1 g151(.A (data_in[5]), .B (n_0), .Y (n_3));
  XNOR2X1 g152(.A (data_in[6]), .B (data_in[5]), .Y (n_2));
  XNOR2X1 g153(.A (data_in[7]), .B (data_in[6]), .Y (n_1));
  XNOR2X1 g154(.A (data_in[4]), .B (data_in[7]), .Y (n_0));
endmodule

module crc_chk_DATA_WIDTH8_POLYNOMIAL_BITS4(clk, rst_n, data_in,
     crc_in, data_out, err_detected, err_corrected);
  input clk, rst_n;
  input [7:0] data_in;
  input [3:0] crc_in;
  output [7:0] data_out;
  output err_detected, err_corrected;
  wire clk, rst_n;
  wire [7:0] data_in;
  wire [3:0] crc_in;
  wire [7:0] data_out;
  wire err_detected, err_corrected;
  wire [3:0] crc_calc;
  wire UNCONNECTED_HIER_Z3, UNCONNECTED_HIER_Z4, n_0, n_1, n_2, n_3,
       n_4, n_5;
  wire n_6;
  crc_gen_DATA_WIDTH8_POLYNOMIAL_BITS4 crc_gen_i(.clk
       (UNCONNECTED_HIER_Z3), .rst_n (UNCONNECTED_HIER_Z4), .data_in
       (data_in), .crc_val (crc_calc));
  DFFRHQX1 err_detected_reg(.RN (rst_n), .CK (clk), .D (n_6), .Q
       (err_detected));
  NAND4XL g134(.A (n_4), .B (n_2), .C (n_5), .D (n_3), .Y (n_6));
  AOI22X1 g135(.A0 (crc_in[0]), .A1 (n_1), .B0 (crc_in[2]), .B1 (n_0),
       .Y (n_5));
  OA22X1 g136(.A0 (crc_in[0]), .A1 (n_1), .B0 (crc_in[2]), .B1 (n_0),
       .Y (n_4));
  XNOR2X1 g137(.A (crc_in[1]), .B (crc_calc[1]), .Y (n_3));
  XNOR2X1 g138(.A (crc_in[3]), .B (crc_calc[3]), .Y (n_2));
  INVX1 g139(.A (crc_calc[0]), .Y (n_1));
  INVX1 g140(.A (crc_calc[2]), .Y (n_0));
endmodule

module crc_gen_DATA_WIDTH8_POLYNOMIAL_BITS4_3(clk, rst_n, data_in,
     crc_val);
  input clk, rst_n;
  input [7:0] data_in;
  output [3:0] crc_val;
  wire clk, rst_n;
  wire [7:0] data_in;
  wire [3:0] crc_val;
  wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_8;
  XNOR2X1 g139(.A (n_6), .B (crc_val[0]), .Y (crc_val[1]));
  XNOR2X1 g140(.A (n_5), .B (n_6), .Y (crc_val[2]));
  CLKXOR2X1 g141(.A (data_in[0]), .B (n_8), .Y (crc_val[0]));
  XNOR2X1 g142(.A (n_0), .B (n_4), .Y (n_8));
  XOR2XL g143(.A (n_4), .B (n_5), .Y (crc_val[3]));
  XNOR2X1 g144(.A (data_in[1]), .B (n_3), .Y (n_6));
  XNOR2X1 g145(.A (data_in[2]), .B (n_2), .Y (n_5));
  XNOR2X1 g146(.A (data_in[3]), .B (n_1), .Y (n_4));
  XNOR2X1 g147(.A (data_in[5]), .B (n_0), .Y (n_3));
  XNOR2X1 g148(.A (data_in[5]), .B (data_in[6]), .Y (n_2));
  XNOR2X1 g149(.A (data_in[6]), .B (data_in[7]), .Y (n_1));
  XNOR2X1 g150(.A (data_in[4]), .B (data_in[7]), .Y (n_0));
endmodule

module mem_with_crc_DATA_WIDTH8_POLYNOMIAL_BITS4(clk, rst_n, mem_wr,
     mem_data_in, crc_data_in, mem_data_out, crc_data_out);
  input clk, rst_n, mem_wr;
  input [7:0] mem_data_in;
  input [3:0] crc_data_in;
  output [7:0] mem_data_out;
  output [3:0] crc_data_out;
  wire clk, rst_n, mem_wr;
  wire [7:0] mem_data_in;
  wire [3:0] crc_data_in;
  wire [7:0] mem_data_out;
  wire [3:0] crc_data_out;
  wire n_0, n_1, n_2, n_3, n_4, n_5, n_6, n_7;
  wire n_8, n_9, n_10, n_11;
  DFFRHQX1 mem_crc_reg_0(.RN (rst_n), .CK (clk), .D (n_10), .Q
       (crc_data_out[0]));
  DFFRHQX1 mem_crc_reg_1(.RN (rst_n), .CK (clk), .D (n_8), .Q
       (crc_data_out[1]));
  DFFRHQX1 mem_reg_4(.RN (rst_n), .CK (clk), .D (n_0), .Q
       (mem_data_out[4]));
  DFFRHQX1 mem_reg_5(.RN (rst_n), .CK (clk), .D (n_11), .Q
       (mem_data_out[5]));
  DFFRHQX1 mem_reg_6(.RN (rst_n), .CK (clk), .D (n_9), .Q
       (mem_data_out[6]));
  DFFRHQX1 mem_reg_7(.RN (rst_n), .CK (clk), .D (n_6), .Q
       (mem_data_out[7]));
  DFFRHQX1 mem_crc_reg_2(.RN (rst_n), .CK (clk), .D (n_7), .Q
       (crc_data_out[2]));
  DFFRHQX1 mem_crc_reg_3(.RN (rst_n), .CK (clk), .D (n_5), .Q
       (crc_data_out[3]));
  DFFRHQX1 mem_reg_0(.RN (rst_n), .CK (clk), .D (n_4), .Q
       (mem_data_out[0]));
  DFFRHQX1 mem_reg_1(.RN (rst_n), .CK (clk), .D (n_3), .Q
       (mem_data_out[1]));
  DFFRHQX1 mem_reg_2(.RN (rst_n), .CK (clk), .D (n_2), .Q
       (mem_data_out[2]));
  DFFRHQX1 mem_reg_3(.RN (rst_n), .CK (clk), .D (n_1), .Q
       (mem_data_out[3]));
  MX2XL g28(.A (mem_data_out[5]), .B (mem_data_in[5]), .S0 (mem_wr), .Y
       (n_11));
  MX2XL g29(.A (crc_data_out[0]), .B (crc_data_in[0]), .S0 (mem_wr), .Y
       (n_10));
  MX2XL g30(.A (mem_data_out[6]), .B (mem_data_in[6]), .S0 (mem_wr), .Y
       (n_9));
  MX2XL g31(.A (crc_data_out[1]), .B (crc_data_in[1]), .S0 (mem_wr), .Y
       (n_8));
  MX2XL g32(.A (crc_data_out[2]), .B (crc_data_in[2]), .S0 (mem_wr), .Y
       (n_7));
  MX2XL g33(.A (mem_data_out[7]), .B (mem_data_in[7]), .S0 (mem_wr), .Y
       (n_6));
  MX2XL g34(.A (crc_data_out[3]), .B (crc_data_in[3]), .S0 (mem_wr), .Y
       (n_5));
  MX2XL g35(.A (mem_data_out[0]), .B (mem_data_in[0]), .S0 (mem_wr), .Y
       (n_4));
  MX2XL g36(.A (mem_data_out[1]), .B (mem_data_in[1]), .S0 (mem_wr), .Y
       (n_3));
  MX2XL g37(.A (mem_data_out[2]), .B (mem_data_in[2]), .S0 (mem_wr), .Y
       (n_2));
  MX2XL g38(.A (mem_data_out[3]), .B (mem_data_in[3]), .S0 (mem_wr), .Y
       (n_1));
  MX2XL g39(.A (mem_data_out[4]), .B (mem_data_in[4]), .S0 (mem_wr), .Y
       (n_0));
endmodule

module crc_mem_DATA_WIDTH8_POLYNOMIAL_BITS4_OUTPUT_FF0(clk, rst_n,
     mem_wr, mem_data_in, mem_data_out, err_detected, err_corrected);
  input clk, rst_n, mem_wr;
  input [7:0] mem_data_in;
  output [7:0] mem_data_out;
  output err_detected, err_corrected;
  wire clk, rst_n, mem_wr;
  wire [7:0] mem_data_in;
  wire [7:0] mem_data_out;
  wire err_detected, err_corrected;
  wire [3:0] mem_crc;
  wire [3:0] crc_wr;
  wire UNCONNECTED32, UNCONNECTED33, UNCONNECTED34, UNCONNECTED35,
       UNCONNECTED36, UNCONNECTED37, UNCONNECTED38, UNCONNECTED39;
  wire UNCONNECTED40, UNCONNECTED_HIER_Z5, UNCONNECTED_HIER_Z6;
  crc_chk_DATA_WIDTH8_POLYNOMIAL_BITS4 crc_chk_i(.clk (clk), .rst_n
       (rst_n), .data_in (mem_data_out), .crc_in (mem_crc), .data_out
       ({UNCONNECTED39, UNCONNECTED38, UNCONNECTED37, UNCONNECTED36,
       UNCONNECTED35, UNCONNECTED34, UNCONNECTED33, UNCONNECTED32}),
       .err_detected (err_detected), .err_corrected (UNCONNECTED40));
  crc_gen_DATA_WIDTH8_POLYNOMIAL_BITS4_3 crc_gen_wr_i(.clk
       (UNCONNECTED_HIER_Z5), .rst_n (UNCONNECTED_HIER_Z6), .data_in
       (mem_data_in), .crc_val (crc_wr));
  mem_with_crc_DATA_WIDTH8_POLYNOMIAL_BITS4 mem_with_crc_i(.clk (clk),
       .rst_n (rst_n), .mem_wr (mem_wr), .mem_data_in (mem_data_in),
       .crc_data_in (crc_wr), .mem_data_out (mem_data_out),
       .crc_data_out (mem_crc));
endmodule

module dut(clk, rst_n, mem1_wr, mem1_data_in, mem1_data_out,
     mem1_err_detected, mem1_err_corrected, mem2_wr, mem2_data_in,
     mem2_data_out, mem2_err_detected, mem2_err_corrected);
  input clk, rst_n, mem1_wr, mem2_wr;
  input [31:0] mem1_data_in;
  input [7:0] mem2_data_in;
  output [31:0] mem1_data_out;
  output mem1_err_detected, mem1_err_corrected, mem2_err_detected,
       mem2_err_corrected;
  output [7:0] mem2_data_out;
  wire clk, rst_n, mem1_wr, mem2_wr;
  wire [31:0] mem1_data_in;
  wire [7:0] mem2_data_in;
  wire [31:0] mem1_data_out;
  wire mem1_err_detected, mem1_err_corrected, mem2_err_detected,
       mem2_err_corrected;
  wire [7:0] mem2_data_out;
  wire UNCONNECTED41, UNCONNECTED42;
  assign mem2_err_corrected = 1'b0;
  assign mem1_err_corrected = 1'b0;
  crc_mem_DATA_WIDTH32_POLYNOMIAL_BITS8_OUTPUT_FF1 mem1_i(.clk (clk),
       .rst_n (rst_n), .mem_wr (mem1_wr), .mem_data_in (mem1_data_in),
       .mem_data_out (mem1_data_out), .err_detected
       (mem1_err_detected), .err_corrected (UNCONNECTED41));
  crc_mem_DATA_WIDTH8_POLYNOMIAL_BITS4_OUTPUT_FF0 mem2_i(.clk (clk),
       .rst_n (rst_n), .mem_wr (mem2_wr), .mem_data_in (mem2_data_in),
       .mem_data_out (mem2_data_out), .err_detected
       (mem2_err_detected), .err_corrected (UNCONNECTED42));
endmodule

