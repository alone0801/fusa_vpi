
//&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&
// GF(5) Error pattern ROM
//&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&&

function[30:0] fn_err_pat_dcd_gf5_rom;						
input[9:0] syndromes; 

reg[30:0] errs;   
begin
 case(syndromes)  

10'h369 : errs =          31'b0000000000000000000000000000001; // S (0x00000001) 
//10'h2d2 : errs =          31'b0000000000000000000000000000011; // D (0x00000003) 
//10'h01f : errs =          31'b0000000000000000000000000000101; // D (0x00000005) 
//10'h2ec : errs =          31'b0000000000000000000000000001001; // D (0x00000009) 
//10'h063 : errs =          31'b0000000000000000000000000010001; // D (0x00000011) 
//10'h214 : errs =          31'b0000000000000000000000000100001; // D (0x00000021) 
//10'h193 : errs =          31'b0000000000000000000000001000001; // D (0x00000041) 
//10'h1f4 : errs =          31'b0000000000000000000000010000001; // D (0x00000081) 
//10'h13a : errs =          31'b0000000000000000000000100000001; // D (0x00000101) 
//10'h0a6 : errs =          31'b0000000000000000000001000000001; // D (0x00000201) 
//10'h39e : errs =          31'b0000000000000000000010000000001; // D (0x00000401) 
//10'h287 : errs =          31'b0000000000000000000100000000001; // D (0x00000801) 
//10'h0b5 : errs =          31'b0000000000000000001000000000001; // D (0x00001001) 
//10'h3b8 : errs =          31'b0000000000000000010000000000001; // D (0x00002001) 
//10'h2cb : errs =          31'b0000000000000000100000000000001; // D (0x00004001) 
//10'h02d : errs =          31'b0000000000000001000000000000001; // D (0x00008001) 
//10'h288 : errs =          31'b0000000000000010000000000000001; // D (0x00010001) 
//10'h0ab : errs =          31'b0000000000000100000000000000001; // D (0x00020001) 
//10'h384 : errs =          31'b0000000000001000000000000000001; // D (0x00040001) 
//10'h2b3 : errs =          31'b0000000000010000000000000000001; // D (0x00080001) 
//10'h0dd : errs =          31'b0000000000100000000000000000001; // D (0x00100001) 
//10'h368 : errs =          31'b0000000001000000000000000000001; // D (0x00200001) 
//10'h36b : errs =          31'b0000000010000000000000000000001; // D (0x00400001) 
//10'h36d : errs =          31'b0000000100000000000000000000001; // D (0x00800001) 
//10'h361 : errs =          31'b0000001000000000000000000000001; // D (0x01000001) 
//10'h379 : errs =          31'b0000010000000000000000000000001; // D (0x02000001) 
//10'h349 : errs =          31'b0000100000000000000000000000001; // D (0x04000001) 
//10'h329 : errs =          31'b0001000000000000000000000000001; // D (0x08000001) 
//10'h3e9 : errs =          31'b0010000000000000000000000000001; // D (0x10000001) 
//10'h269 : errs =          31'b0100000000000000000000000000001; // D (0x20000001) 
//10'h169 : errs =          31'b1000000000000000000000000000001; // D (0x40000001) 
10'h2d2 : errs =          31'b0000000000000000000000000000011; // D (0x00000003) 
10'h1bb : errs =          31'b0000000000000000000000000000010; // S (0x00000002) 
//10'h2cd : errs =          31'b0000000000000000000000000000110; // D (0x00000006) 
//10'h03e : errs =          31'b0000000000000000000000000001010; // D (0x0000000a) 
//10'h2b1 : errs =          31'b0000000000000000000000000010010; // D (0x00000012) 
//10'h0c6 : errs =          31'b0000000000000000000000000100010; // D (0x00000022) 
//10'h341 : errs =          31'b0000000000000000000000001000010; // D (0x00000042) 
//10'h326 : errs =          31'b0000000000000000000000010000010; // D (0x00000082) 
//10'h3e8 : errs =          31'b0000000000000000000000100000010; // D (0x00000102) 
//10'h274 : errs =          31'b0000000000000000000001000000010; // D (0x00000202) 
//10'h14c : errs =          31'b0000000000000000000010000000010; // D (0x00000402) 
//10'h055 : errs =          31'b0000000000000000000100000000010; // D (0x00000802) 
//10'h267 : errs =          31'b0000000000000000001000000000010; // D (0x00001002) 
//10'h16a : errs =          31'b0000000000000000010000000000010; // D (0x00002002) 
//10'h019 : errs =          31'b0000000000000000100000000000010; // D (0x00004002) 
//10'h2ff : errs =          31'b0000000000000001000000000000010; // D (0x00008002) 
//10'h05a : errs =          31'b0000000000000010000000000000010; // D (0x00010002) 
//10'h279 : errs =          31'b0000000000000100000000000000010; // D (0x00020002) 
//10'h156 : errs =          31'b0000000000001000000000000000010; // D (0x00040002) 
//10'h061 : errs =          31'b0000000000010000000000000000010; // D (0x00080002) 
//10'h20f : errs =          31'b0000000000100000000000000000010; // D (0x00100002) 
//10'h1ba : errs =          31'b0000000001000000000000000000010; // D (0x00200002) 
//10'h1b9 : errs =          31'b0000000010000000000000000000010; // D (0x00400002) 
//10'h1bf : errs =          31'b0000000100000000000000000000010; // D (0x00800002) 
//10'h1b3 : errs =          31'b0000001000000000000000000000010; // D (0x01000002) 
//10'h1ab : errs =          31'b0000010000000000000000000000010; // D (0x02000002) 
//10'h19b : errs =          31'b0000100000000000000000000000010; // D (0x04000002) 
//10'h1fb : errs =          31'b0001000000000000000000000000010; // D (0x08000002) 
//10'h13b : errs =          31'b0010000000000000000000000000010; // D (0x10000002) 
//10'h0bb : errs =          31'b0100000000000000000000000000010; // D (0x20000002) 
//10'h3bb : errs =          31'b1000000000000000000000000000010; // D (0x40000002) 
10'h01f : errs =          31'b0000000000000000000000000000101; // D (0x00000005) 
10'h2cd : errs =          31'b0000000000000000000000000000110; // D (0x00000006) 
10'h376 : errs =          31'b0000000000000000000000000000100; // S (0x00000004) 
//10'h2f3 : errs =          31'b0000000000000000000000000001100; // D (0x0000000c) 
//10'h07c : errs =          31'b0000000000000000000000000010100; // D (0x00000014) 
//10'h20b : errs =          31'b0000000000000000000000000100100; // D (0x00000024) 
//10'h18c : errs =          31'b0000000000000000000000001000100; // D (0x00000044) 
//10'h1eb : errs =          31'b0000000000000000000000010000100; // D (0x00000084) 
//10'h125 : errs =          31'b0000000000000000000000100000100; // D (0x00000104) 
//10'h0b9 : errs =          31'b0000000000000000000001000000100; // D (0x00000204) 
//10'h381 : errs =          31'b0000000000000000000010000000100; // D (0x00000404) 
//10'h298 : errs =          31'b0000000000000000000100000000100; // D (0x00000804) 
//10'h0aa : errs =          31'b0000000000000000001000000000100; // D (0x00001004) 
//10'h3a7 : errs =          31'b0000000000000000010000000000100; // D (0x00002004) 
//10'h2d4 : errs =          31'b0000000000000000100000000000100; // D (0x00004004) 
//10'h032 : errs =          31'b0000000000000001000000000000100; // D (0x00008004) 
//10'h297 : errs =          31'b0000000000000010000000000000100; // D (0x00010004) 
//10'h0b4 : errs =          31'b0000000000000100000000000000100; // D (0x00020004) 
//10'h39b : errs =          31'b0000000000001000000000000000100; // D (0x00040004) 
//10'h2ac : errs =          31'b0000000000010000000000000000100; // D (0x00080004) 
//10'h0c2 : errs =          31'b0000000000100000000000000000100; // D (0x00100004) 
//10'h377 : errs =          31'b0000000001000000000000000000100; // D (0x00200004) 
//10'h374 : errs =          31'b0000000010000000000000000000100; // D (0x00400004) 
//10'h372 : errs =          31'b0000000100000000000000000000100; // D (0x00800004) 
//10'h37e : errs =          31'b0000001000000000000000000000100; // D (0x01000004) 
//10'h366 : errs =          31'b0000010000000000000000000000100; // D (0x02000004) 
//10'h356 : errs =          31'b0000100000000000000000000000100; // D (0x04000004) 
//10'h336 : errs =          31'b0001000000000000000000000000100; // D (0x08000004) 
//10'h3f6 : errs =          31'b0010000000000000000000000000100; // D (0x10000004) 
//10'h276 : errs =          31'b0100000000000000000000000000100; // D (0x20000004) 
//10'h176 : errs =          31'b1000000000000000000000000000100; // D (0x40000004) 
10'h2ec : errs =          31'b0000000000000000000000000001001; // D (0x00000009) 
10'h03e : errs =          31'b0000000000000000000000000001010; // D (0x0000000a) 
10'h2f3 : errs =          31'b0000000000000000000000000001100; // D (0x0000000c) 
10'h185 : errs =          31'b0000000000000000000000000001000; // S (0x00000008) 
//10'h28f : errs =          31'b0000000000000000000000000011000; // D (0x00000018) 
//10'h0f8 : errs =          31'b0000000000000000000000000101000; // D (0x00000028) 
//10'h37f : errs =          31'b0000000000000000000000001001000; // D (0x00000048) 
//10'h318 : errs =          31'b0000000000000000000000010001000; // D (0x00000088) 
//10'h3d6 : errs =          31'b0000000000000000000000100001000; // D (0x00000108) 
//10'h24a : errs =          31'b0000000000000000000001000001000; // D (0x00000208) 
//10'h172 : errs =          31'b0000000000000000000010000001000; // D (0x00000408) 
//10'h06b : errs =          31'b0000000000000000000100000001000; // D (0x00000808) 
//10'h259 : errs =          31'b0000000000000000001000000001000; // D (0x00001008) 
//10'h154 : errs =          31'b0000000000000000010000000001000; // D (0x00002008) 
//10'h027 : errs =          31'b0000000000000000100000000001000; // D (0x00004008) 
//10'h2c1 : errs =          31'b0000000000000001000000000001000; // D (0x00008008) 
//10'h064 : errs =          31'b0000000000000010000000000001000; // D (0x00010008) 
//10'h247 : errs =          31'b0000000000000100000000000001000; // D (0x00020008) 
//10'h168 : errs =          31'b0000000000001000000000000001000; // D (0x00040008) 
//10'h05f : errs =          31'b0000000000010000000000000001000; // D (0x00080008) 
//10'h231 : errs =          31'b0000000000100000000000000001000; // D (0x00100008) 
//10'h184 : errs =          31'b0000000001000000000000000001000; // D (0x00200008) 
//10'h187 : errs =          31'b0000000010000000000000000001000; // D (0x00400008) 
//10'h181 : errs =          31'b0000000100000000000000000001000; // D (0x00800008) 
//10'h18d : errs =          31'b0000001000000000000000000001000; // D (0x01000008) 
//10'h195 : errs =          31'b0000010000000000000000000001000; // D (0x02000008) 
//10'h1a5 : errs =          31'b0000100000000000000000000001000; // D (0x04000008) 
//10'h1c5 : errs =          31'b0001000000000000000000000001000; // D (0x08000008) 
//10'h105 : errs =          31'b0010000000000000000000000001000; // D (0x10000008) 
//10'h085 : errs =          31'b0100000000000000000000000001000; // D (0x20000008) 
//10'h385 : errs =          31'b1000000000000000000000000001000; // D (0x40000008) 
10'h063 : errs =          31'b0000000000000000000000000010001; // D (0x00000011) 
10'h2b1 : errs =          31'b0000000000000000000000000010010; // D (0x00000012) 
10'h07c : errs =          31'b0000000000000000000000000010100; // D (0x00000014) 
10'h28f : errs =          31'b0000000000000000000000000011000; // D (0x00000018) 
10'h30a : errs =          31'b0000000000000000000000000010000; // S (0x00000010) 
//10'h277 : errs =          31'b0000000000000000000000000110000; // D (0x00000030) 
//10'h1f0 : errs =          31'b0000000000000000000000001010000; // D (0x00000050) 
//10'h197 : errs =          31'b0000000000000000000000010010000; // D (0x00000090) 
//10'h159 : errs =          31'b0000000000000000000000100010000; // D (0x00000110) 
//10'h0c5 : errs =          31'b0000000000000000000001000010000; // D (0x00000210) 
//10'h3fd : errs =          31'b0000000000000000000010000010000; // D (0x00000410) 
//10'h2e4 : errs =          31'b0000000000000000000100000010000; // D (0x00000810) 
//10'h0d6 : errs =          31'b0000000000000000001000000010000; // D (0x00001010) 
//10'h3db : errs =          31'b0000000000000000010000000010000; // D (0x00002010) 
//10'h2a8 : errs =          31'b0000000000000000100000000010000; // D (0x00004010) 
//10'h04e : errs =          31'b0000000000000001000000000010000; // D (0x00008010) 
//10'h2eb : errs =          31'b0000000000000010000000000010000; // D (0x00010010) 
//10'h0c8 : errs =          31'b0000000000000100000000000010000; // D (0x00020010) 
//10'h3e7 : errs =          31'b0000000000001000000000000010000; // D (0x00040010) 
//10'h2d0 : errs =          31'b0000000000010000000000000010000; // D (0x00080010) 
//10'h0be : errs =          31'b0000000000100000000000000010000; // D (0x00100010) 
//10'h30b : errs =          31'b0000000001000000000000000010000; // D (0x00200010) 
//10'h308 : errs =          31'b0000000010000000000000000010000; // D (0x00400010) 
//10'h30e : errs =          31'b0000000100000000000000000010000; // D (0x00800010) 
//10'h302 : errs =          31'b0000001000000000000000000010000; // D (0x01000010) 
//10'h31a : errs =          31'b0000010000000000000000000010000; // D (0x02000010) 
//10'h32a : errs =          31'b0000100000000000000000000010000; // D (0x04000010) 
//10'h34a : errs =          31'b0001000000000000000000000010000; // D (0x08000010) 
//10'h38a : errs =          31'b0010000000000000000000000010000; // D (0x10000010) 
//10'h20a : errs =          31'b0100000000000000000000000010000; // D (0x20000010) 
//10'h10a : errs =          31'b1000000000000000000000000010000; // D (0x40000010) 
10'h214 : errs =          31'b0000000000000000000000000100001; // D (0x00000021) 
10'h0c6 : errs =          31'b0000000000000000000000000100010; // D (0x00000022) 
10'h20b : errs =          31'b0000000000000000000000000100100; // D (0x00000024) 
10'h0f8 : errs =          31'b0000000000000000000000000101000; // D (0x00000028) 
10'h277 : errs =          31'b0000000000000000000000000110000; // D (0x00000030) 
10'h17d : errs =          31'b0000000000000000000000000100000; // S (0x00000020) 
//10'h387 : errs =          31'b0000000000000000000000001100000; // D (0x00000060) 
//10'h3e0 : errs =          31'b0000000000000000000000010100000; // D (0x000000a0) 
//10'h32e : errs =          31'b0000000000000000000000100100000; // D (0x00000120) 
//10'h2b2 : errs =          31'b0000000000000000000001000100000; // D (0x00000220) 
//10'h18a : errs =          31'b0000000000000000000010000100000; // D (0x00000420) 
//10'h093 : errs =          31'b0000000000000000000100000100000; // D (0x00000820) 
//10'h2a1 : errs =          31'b0000000000000000001000000100000; // D (0x00001020) 
//10'h1ac : errs =          31'b0000000000000000010000000100000; // D (0x00002020) 
//10'h0df : errs =          31'b0000000000000000100000000100000; // D (0x00004020) 
//10'h239 : errs =          31'b0000000000000001000000000100000; // D (0x00008020) 
//10'h09c : errs =          31'b0000000000000010000000000100000; // D (0x00010020) 
//10'h2bf : errs =          31'b0000000000000100000000000100000; // D (0x00020020) 
//10'h190 : errs =          31'b0000000000001000000000000100000; // D (0x00040020) 
//10'h0a7 : errs =          31'b0000000000010000000000000100000; // D (0x00080020) 
//10'h2c9 : errs =          31'b0000000000100000000000000100000; // D (0x00100020) 
//10'h17c : errs =          31'b0000000001000000000000000100000; // D (0x00200020) 
//10'h17f : errs =          31'b0000000010000000000000000100000; // D (0x00400020) 
//10'h179 : errs =          31'b0000000100000000000000000100000; // D (0x00800020) 
//10'h175 : errs =          31'b0000001000000000000000000100000; // D (0x01000020) 
//10'h16d : errs =          31'b0000010000000000000000000100000; // D (0x02000020) 
//10'h15d : errs =          31'b0000100000000000000000000100000; // D (0x04000020) 
//10'h13d : errs =          31'b0001000000000000000000000100000; // D (0x08000020) 
//10'h1fd : errs =          31'b0010000000000000000000000100000; // D (0x10000020) 
//10'h07d : errs =          31'b0100000000000000000000000100000; // D (0x20000020) 
//10'h37d : errs =          31'b1000000000000000000000000100000; // D (0x40000020) 
10'h193 : errs =          31'b0000000000000000000000001000001; // D (0x00000041) 
10'h341 : errs =          31'b0000000000000000000000001000010; // D (0x00000042) 
10'h18c : errs =          31'b0000000000000000000000001000100; // D (0x00000044) 
10'h37f : errs =          31'b0000000000000000000000001001000; // D (0x00000048) 
10'h1f0 : errs =          31'b0000000000000000000000001010000; // D (0x00000050) 
10'h387 : errs =          31'b0000000000000000000000001100000; // D (0x00000060) 
10'h2fa : errs =          31'b0000000000000000000000001000000; // S (0x00000040) 
//10'h067 : errs =          31'b0000000000000000000000011000000; // D (0x000000c0) 
//10'h0a9 : errs =          31'b0000000000000000000000101000000; // D (0x00000140) 
//10'h135 : errs =          31'b0000000000000000000001001000000; // D (0x00000240) 
//10'h20d : errs =          31'b0000000000000000000010001000000; // D (0x00000440) 
//10'h314 : errs =          31'b0000000000000000000100001000000; // D (0x00000840) 
//10'h126 : errs =          31'b0000000000000000001000001000000; // D (0x00001040) 
//10'h22b : errs =          31'b0000000000000000010000001000000; // D (0x00002040) 
//10'h358 : errs =          31'b0000000000000000100000001000000; // D (0x00004040) 
//10'h1be : errs =          31'b0000000000000001000000001000000; // D (0x00008040) 
//10'h31b : errs =          31'b0000000000000010000000001000000; // D (0x00010040) 
//10'h138 : errs =          31'b0000000000000100000000001000000; // D (0x00020040) 
//10'h217 : errs =          31'b0000000000001000000000001000000; // D (0x00040040) 
//10'h320 : errs =          31'b0000000000010000000000001000000; // D (0x00080040) 
//10'h14e : errs =          31'b0000000000100000000000001000000; // D (0x00100040) 
//10'h2fb : errs =          31'b0000000001000000000000001000000; // D (0x00200040) 
//10'h2f8 : errs =          31'b0000000010000000000000001000000; // D (0x00400040) 
//10'h2fe : errs =          31'b0000000100000000000000001000000; // D (0x00800040) 
//10'h2f2 : errs =          31'b0000001000000000000000001000000; // D (0x01000040) 
//10'h2ea : errs =          31'b0000010000000000000000001000000; // D (0x02000040) 
//10'h2da : errs =          31'b0000100000000000000000001000000; // D (0x04000040) 
//10'h2ba : errs =          31'b0001000000000000000000001000000; // D (0x08000040) 
//10'h27a : errs =          31'b0010000000000000000000001000000; // D (0x10000040) 
//10'h3fa : errs =          31'b0100000000000000000000001000000; // D (0x20000040) 
//10'h0fa : errs =          31'b1000000000000000000000001000000; // D (0x40000040) 
10'h1f4 : errs =          31'b0000000000000000000000010000001; // D (0x00000081) 
10'h326 : errs =          31'b0000000000000000000000010000010; // D (0x00000082) 
10'h1eb : errs =          31'b0000000000000000000000010000100; // D (0x00000084) 
10'h318 : errs =          31'b0000000000000000000000010001000; // D (0x00000088) 
10'h197 : errs =          31'b0000000000000000000000010010000; // D (0x00000090) 
10'h3e0 : errs =          31'b0000000000000000000000010100000; // D (0x000000a0) 
10'h067 : errs =          31'b0000000000000000000000011000000; // D (0x000000c0) 
10'h29d : errs =          31'b0000000000000000000000010000000; // S (0x00000080) 
//10'h0ce : errs =          31'b0000000000000000000000110000000; // D (0x00000180) 
//10'h152 : errs =          31'b0000000000000000000001010000000; // D (0x00000280) 
//10'h26a : errs =          31'b0000000000000000000010010000000; // D (0x00000480) 
//10'h373 : errs =          31'b0000000000000000000100010000000; // D (0x00000880) 
//10'h141 : errs =          31'b0000000000000000001000010000000; // D (0x00001080) 
//10'h24c : errs =          31'b0000000000000000010000010000000; // D (0x00002080) 
//10'h33f : errs =          31'b0000000000000000100000010000000; // D (0x00004080) 
//10'h1d9 : errs =          31'b0000000000000001000000010000000; // D (0x00008080) 
//10'h37c : errs =          31'b0000000000000010000000010000000; // D (0x00010080) 
//10'h15f : errs =          31'b0000000000000100000000010000000; // D (0x00020080) 
//10'h270 : errs =          31'b0000000000001000000000010000000; // D (0x00040080) 
//10'h347 : errs =          31'b0000000000010000000000010000000; // D (0x00080080) 
//10'h129 : errs =          31'b0000000000100000000000010000000; // D (0x00100080) 
//10'h29c : errs =          31'b0000000001000000000000010000000; // D (0x00200080) 
//10'h29f : errs =          31'b0000000010000000000000010000000; // D (0x00400080) 
//10'h299 : errs =          31'b0000000100000000000000010000000; // D (0x00800080) 
//10'h295 : errs =          31'b0000001000000000000000010000000; // D (0x01000080) 
//10'h28d : errs =          31'b0000010000000000000000010000000; // D (0x02000080) 
//10'h2bd : errs =          31'b0000100000000000000000010000000; // D (0x04000080) 
//10'h2dd : errs =          31'b0001000000000000000000010000000; // D (0x08000080) 
//10'h21d : errs =          31'b0010000000000000000000010000000; // D (0x10000080) 
//10'h39d : errs =          31'b0100000000000000000000010000000; // D (0x20000080) 
//10'h09d : errs =          31'b1000000000000000000000010000000; // D (0x40000080) 
10'h13a : errs =          31'b0000000000000000000000100000001; // D (0x00000101) 
10'h3e8 : errs =          31'b0000000000000000000000100000010; // D (0x00000102) 
10'h125 : errs =          31'b0000000000000000000000100000100; // D (0x00000104) 
10'h3d6 : errs =          31'b0000000000000000000000100001000; // D (0x00000108) 
10'h159 : errs =          31'b0000000000000000000000100010000; // D (0x00000110) 
10'h32e : errs =          31'b0000000000000000000000100100000; // D (0x00000120) 
10'h0a9 : errs =          31'b0000000000000000000000101000000; // D (0x00000140) 
10'h0ce : errs =          31'b0000000000000000000000110000000; // D (0x00000180) 
10'h253 : errs =          31'b0000000000000000000000100000000; // S (0x00000100) 
//10'h19c : errs =          31'b0000000000000000000001100000000; // D (0x00000300) 
//10'h2a4 : errs =          31'b0000000000000000000010100000000; // D (0x00000500) 
//10'h3bd : errs =          31'b0000000000000000000100100000000; // D (0x00000900) 
//10'h18f : errs =          31'b0000000000000000001000100000000; // D (0x00001100) 
//10'h282 : errs =          31'b0000000000000000010000100000000; // D (0x00002100) 
//10'h3f1 : errs =          31'b0000000000000000100000100000000; // D (0x00004100) 
//10'h117 : errs =          31'b0000000000000001000000100000000; // D (0x00008100) 
//10'h3b2 : errs =          31'b0000000000000010000000100000000; // D (0x00010100) 
//10'h191 : errs =          31'b0000000000000100000000100000000; // D (0x00020100) 
//10'h2be : errs =          31'b0000000000001000000000100000000; // D (0x00040100) 
//10'h389 : errs =          31'b0000000000010000000000100000000; // D (0x00080100) 
//10'h1e7 : errs =          31'b0000000000100000000000100000000; // D (0x00100100) 
//10'h252 : errs =          31'b0000000001000000000000100000000; // D (0x00200100) 
//10'h251 : errs =          31'b0000000010000000000000100000000; // D (0x00400100) 
//10'h257 : errs =          31'b0000000100000000000000100000000; // D (0x00800100) 
//10'h25b : errs =          31'b0000001000000000000000100000000; // D (0x01000100) 
//10'h243 : errs =          31'b0000010000000000000000100000000; // D (0x02000100) 
//10'h273 : errs =          31'b0000100000000000000000100000000; // D (0x04000100) 
//10'h213 : errs =          31'b0001000000000000000000100000000; // D (0x08000100) 
//10'h2d3 : errs =          31'b0010000000000000000000100000000; // D (0x10000100) 
//10'h353 : errs =          31'b0100000000000000000000100000000; // D (0x20000100) 
//10'h053 : errs =          31'b1000000000000000000000100000000; // D (0x40000100) 
10'h0a6 : errs =          31'b0000000000000000000001000000001; // D (0x00000201) 
10'h274 : errs =          31'b0000000000000000000001000000010; // D (0x00000202) 
10'h0b9 : errs =          31'b0000000000000000000001000000100; // D (0x00000204) 
10'h24a : errs =          31'b0000000000000000000001000001000; // D (0x00000208) 
10'h0c5 : errs =          31'b0000000000000000000001000010000; // D (0x00000210) 
10'h2b2 : errs =          31'b0000000000000000000001000100000; // D (0x00000220) 
10'h135 : errs =          31'b0000000000000000000001001000000; // D (0x00000240) 
10'h152 : errs =          31'b0000000000000000000001010000000; // D (0x00000280) 
10'h19c : errs =          31'b0000000000000000000001100000000; // D (0x00000300) 
10'h3cf : errs =          31'b0000000000000000000001000000000; // S (0x00000200) 
//10'h338 : errs =          31'b0000000000000000000011000000000; // D (0x00000600) 
//10'h221 : errs =          31'b0000000000000000000101000000000; // D (0x00000a00) 
//10'h013 : errs =          31'b0000000000000000001001000000000; // D (0x00001200) 
//10'h31e : errs =          31'b0000000000000000010001000000000; // D (0x00002200) 
//10'h26d : errs =          31'b0000000000000000100001000000000; // D (0x00004200) 
//10'h08b : errs =          31'b0000000000000001000001000000000; // D (0x00008200) 
//10'h22e : errs =          31'b0000000000000010000001000000000; // D (0x00010200) 
//10'h00d : errs =          31'b0000000000000100000001000000000; // D (0x00020200) 
//10'h322 : errs =          31'b0000000000001000000001000000000; // D (0x00040200) 
//10'h215 : errs =          31'b0000000000010000000001000000000; // D (0x00080200) 
//10'h07b : errs =          31'b0000000000100000000001000000000; // D (0x00100200) 
//10'h3ce : errs =          31'b0000000001000000000001000000000; // D (0x00200200) 
//10'h3cd : errs =          31'b0000000010000000000001000000000; // D (0x00400200) 
//10'h3cb : errs =          31'b0000000100000000000001000000000; // D (0x00800200) 
//10'h3c7 : errs =          31'b0000001000000000000001000000000; // D (0x01000200) 
//10'h3df : errs =          31'b0000010000000000000001000000000; // D (0x02000200) 
//10'h3ef : errs =          31'b0000100000000000000001000000000; // D (0x04000200) 
//10'h38f : errs =          31'b0001000000000000000001000000000; // D (0x08000200) 
//10'h34f : errs =          31'b0010000000000000000001000000000; // D (0x10000200) 
//10'h2cf : errs =          31'b0100000000000000000001000000000; // D (0x20000200) 
//10'h1cf : errs =          31'b1000000000000000000001000000000; // D (0x40000200) 
10'h39e : errs =          31'b0000000000000000000010000000001; // D (0x00000401) 
10'h14c : errs =          31'b0000000000000000000010000000010; // D (0x00000402) 
10'h381 : errs =          31'b0000000000000000000010000000100; // D (0x00000404) 
10'h172 : errs =          31'b0000000000000000000010000001000; // D (0x00000408) 
10'h3fd : errs =          31'b0000000000000000000010000010000; // D (0x00000410) 
10'h18a : errs =          31'b0000000000000000000010000100000; // D (0x00000420) 
10'h20d : errs =          31'b0000000000000000000010001000000; // D (0x00000440) 
10'h26a : errs =          31'b0000000000000000000010010000000; // D (0x00000480) 
10'h2a4 : errs =          31'b0000000000000000000010100000000; // D (0x00000500) 
10'h338 : errs =          31'b0000000000000000000011000000000; // D (0x00000600) 
10'h0f7 : errs =          31'b0000000000000000000010000000000; // S (0x00000400) 
//10'h119 : errs =          31'b0000000000000000000110000000000; // D (0x00000c00) 
//10'h32b : errs =          31'b0000000000000000001010000000000; // D (0x00001400) 
//10'h026 : errs =          31'b0000000000000000010010000000000; // D (0x00002400) 
//10'h155 : errs =          31'b0000000000000000100010000000000; // D (0x00004400) 
//10'h3b3 : errs =          31'b0000000000000001000010000000000; // D (0x00008400) 
//10'h116 : errs =          31'b0000000000000010000010000000000; // D (0x00010400) 
//10'h335 : errs =          31'b0000000000000100000010000000000; // D (0x00020400) 
//10'h01a : errs =          31'b0000000000001000000010000000000; // D (0x00040400) 
//10'h12d : errs =          31'b0000000000010000000010000000000; // D (0x00080400) 
//10'h343 : errs =          31'b0000000000100000000010000000000; // D (0x00100400) 
//10'h0f6 : errs =          31'b0000000001000000000010000000000; // D (0x00200400) 
//10'h0f5 : errs =          31'b0000000010000000000010000000000; // D (0x00400400) 
//10'h0f3 : errs =          31'b0000000100000000000010000000000; // D (0x00800400) 
//10'h0ff : errs =          31'b0000001000000000000010000000000; // D (0x01000400) 
//10'h0e7 : errs =          31'b0000010000000000000010000000000; // D (0x02000400) 
//10'h0d7 : errs =          31'b0000100000000000000010000000000; // D (0x04000400) 
//10'h0b7 : errs =          31'b0001000000000000000010000000000; // D (0x08000400) 
//10'h077 : errs =          31'b0010000000000000000010000000000; // D (0x10000400) 
//10'h1f7 : errs =          31'b0100000000000000000010000000000; // D (0x20000400) 
//10'h2f7 : errs =          31'b1000000000000000000010000000000; // D (0x40000400) 
10'h287 : errs =          31'b0000000000000000000100000000001; // D (0x00000801) 
10'h055 : errs =          31'b0000000000000000000100000000010; // D (0x00000802) 
10'h298 : errs =          31'b0000000000000000000100000000100; // D (0x00000804) 
10'h06b : errs =          31'b0000000000000000000100000001000; // D (0x00000808) 
10'h2e4 : errs =          31'b0000000000000000000100000010000; // D (0x00000810) 
10'h093 : errs =          31'b0000000000000000000100000100000; // D (0x00000820) 
10'h314 : errs =          31'b0000000000000000000100001000000; // D (0x00000840) 
10'h373 : errs =          31'b0000000000000000000100010000000; // D (0x00000880) 
10'h3bd : errs =          31'b0000000000000000000100100000000; // D (0x00000900) 
10'h221 : errs =          31'b0000000000000000000101000000000; // D (0x00000a00) 
10'h119 : errs =          31'b0000000000000000000110000000000; // D (0x00000c00) 
10'h1ee : errs =          31'b0000000000000000000100000000000; // S (0x00000800) 
//10'h232 : errs =          31'b0000000000000000001100000000000; // D (0x00001800) 
//10'h13f : errs =          31'b0000000000000000010100000000000; // D (0x00002800) 
//10'h04c : errs =          31'b0000000000000000100100000000000; // D (0x00004800) 
//10'h2aa : errs =          31'b0000000000000001000100000000000; // D (0x00008800) 
//10'h00f : errs =          31'b0000000000000010000100000000000; // D (0x00010800) 
//10'h22c : errs =          31'b0000000000000100000100000000000; // D (0x00020800) 
//10'h103 : errs =          31'b0000000000001000000100000000000; // D (0x00040800) 
//10'h034 : errs =          31'b0000000000010000000100000000000; // D (0x00080800) 
//10'h25a : errs =          31'b0000000000100000000100000000000; // D (0x00100800) 
//10'h1ef : errs =          31'b0000000001000000000100000000000; // D (0x00200800) 
//10'h1ec : errs =          31'b0000000010000000000100000000000; // D (0x00400800) 
//10'h1ea : errs =          31'b0000000100000000000100000000000; // D (0x00800800) 
//10'h1e6 : errs =          31'b0000001000000000000100000000000; // D (0x01000800) 
//10'h1fe : errs =          31'b0000010000000000000100000000000; // D (0x02000800) 
//10'h1ce : errs =          31'b0000100000000000000100000000000; // D (0x04000800) 
//10'h1ae : errs =          31'b0001000000000000000100000000000; // D (0x08000800) 
//10'h16e : errs =          31'b0010000000000000000100000000000; // D (0x10000800) 
//10'h0ee : errs =          31'b0100000000000000000100000000000; // D (0x20000800) 
//10'h3ee : errs =          31'b1000000000000000000100000000000; // D (0x40000800) 
10'h0b5 : errs =          31'b0000000000000000001000000000001; // D (0x00001001) 
10'h267 : errs =          31'b0000000000000000001000000000010; // D (0x00001002) 
10'h0aa : errs =          31'b0000000000000000001000000000100; // D (0x00001004) 
10'h259 : errs =          31'b0000000000000000001000000001000; // D (0x00001008) 
10'h0d6 : errs =          31'b0000000000000000001000000010000; // D (0x00001010) 
10'h2a1 : errs =          31'b0000000000000000001000000100000; // D (0x00001020) 
10'h126 : errs =          31'b0000000000000000001000001000000; // D (0x00001040) 
10'h141 : errs =          31'b0000000000000000001000010000000; // D (0x00001080) 
10'h18f : errs =          31'b0000000000000000001000100000000; // D (0x00001100) 
10'h013 : errs =          31'b0000000000000000001001000000000; // D (0x00001200) 
10'h32b : errs =          31'b0000000000000000001010000000000; // D (0x00001400) 
10'h232 : errs =          31'b0000000000000000001100000000000; // D (0x00001800) 
10'h3dc : errs =          31'b0000000000000000001000000000000; // S (0x00001000) 
//10'h30d : errs =          31'b0000000000000000011000000000000; // D (0x00003000) 
//10'h27e : errs =          31'b0000000000000000101000000000000; // D (0x00005000) 
//10'h098 : errs =          31'b0000000000000001001000000000000; // D (0x00009000) 
//10'h23d : errs =          31'b0000000000000010001000000000000; // D (0x00011000) 
//10'h01e : errs =          31'b0000000000000100001000000000000; // D (0x00021000) 
//10'h331 : errs =          31'b0000000000001000001000000000000; // D (0x00041000) 
//10'h206 : errs =          31'b0000000000010000001000000000000; // D (0x00081000) 
//10'h068 : errs =          31'b0000000000100000001000000000000; // D (0x00101000) 
//10'h3dd : errs =          31'b0000000001000000001000000000000; // D (0x00201000) 
//10'h3de : errs =          31'b0000000010000000001000000000000; // D (0x00401000) 
//10'h3d8 : errs =          31'b0000000100000000001000000000000; // D (0x00801000) 
//10'h3d4 : errs =          31'b0000001000000000001000000000000; // D (0x01001000) 
//10'h3cc : errs =          31'b0000010000000000001000000000000; // D (0x02001000) 
//10'h3fc : errs =          31'b0000100000000000001000000000000; // D (0x04001000) 
//10'h39c : errs =          31'b0001000000000000001000000000000; // D (0x08001000) 
//10'h35c : errs =          31'b0010000000000000001000000000000; // D (0x10001000) 
//10'h2dc : errs =          31'b0100000000000000001000000000000; // D (0x20001000) 
//10'h1dc : errs =          31'b1000000000000000001000000000000; // D (0x40001000) 
10'h3b8 : errs =          31'b0000000000000000010000000000001; // D (0x00002001) 
10'h16a : errs =          31'b0000000000000000010000000000010; // D (0x00002002) 
10'h3a7 : errs =          31'b0000000000000000010000000000100; // D (0x00002004) 
10'h154 : errs =          31'b0000000000000000010000000001000; // D (0x00002008) 
10'h3db : errs =          31'b0000000000000000010000000010000; // D (0x00002010) 
10'h1ac : errs =          31'b0000000000000000010000000100000; // D (0x00002020) 
10'h22b : errs =          31'b0000000000000000010000001000000; // D (0x00002040) 
10'h24c : errs =          31'b0000000000000000010000010000000; // D (0x00002080) 
10'h282 : errs =          31'b0000000000000000010000100000000; // D (0x00002100) 
10'h31e : errs =          31'b0000000000000000010001000000000; // D (0x00002200) 
10'h026 : errs =          31'b0000000000000000010010000000000; // D (0x00002400) 
10'h13f : errs =          31'b0000000000000000010100000000000; // D (0x00002800) 
10'h30d : errs =          31'b0000000000000000011000000000000; // D (0x00003000) 
10'h0d1 : errs =          31'b0000000000000000010000000000000; // S (0x00002000) 
//10'h173 : errs =          31'b0000000000000000110000000000000; // D (0x00006000) 
//10'h395 : errs =          31'b0000000000000001010000000000000; // D (0x0000a000) 
//10'h130 : errs =          31'b0000000000000010010000000000000; // D (0x00012000) 
//10'h313 : errs =          31'b0000000000000100010000000000000; // D (0x00022000) 
//10'h03c : errs =          31'b0000000000001000010000000000000; // D (0x00042000) 
//10'h10b : errs =          31'b0000000000010000010000000000000; // D (0x00082000) 
//10'h365 : errs =          31'b0000000000100000010000000000000; // D (0x00102000) 
//10'h0d0 : errs =          31'b0000000001000000010000000000000; // D (0x00202000) 
//10'h0d3 : errs =          31'b0000000010000000010000000000000; // D (0x00402000) 
//10'h0d5 : errs =          31'b0000000100000000010000000000000; // D (0x00802000) 
//10'h0d9 : errs =          31'b0000001000000000010000000000000; // D (0x01002000) 
//10'h0c1 : errs =          31'b0000010000000000010000000000000; // D (0x02002000) 
//10'h0f1 : errs =          31'b0000100000000000010000000000000; // D (0x04002000) 
//10'h091 : errs =          31'b0001000000000000010000000000000; // D (0x08002000) 
//10'h051 : errs =          31'b0010000000000000010000000000000; // D (0x10002000) 
//10'h1d1 : errs =          31'b0100000000000000010000000000000; // D (0x20002000) 
//10'h2d1 : errs =          31'b1000000000000000010000000000000; // D (0x40002000) 
10'h2cb : errs =          31'b0000000000000000100000000000001; // D (0x00004001) 
10'h019 : errs =          31'b0000000000000000100000000000010; // D (0x00004002) 
10'h2d4 : errs =          31'b0000000000000000100000000000100; // D (0x00004004) 
10'h027 : errs =          31'b0000000000000000100000000001000; // D (0x00004008) 
10'h2a8 : errs =          31'b0000000000000000100000000010000; // D (0x00004010) 
10'h0df : errs =          31'b0000000000000000100000000100000; // D (0x00004020) 
10'h358 : errs =          31'b0000000000000000100000001000000; // D (0x00004040) 
10'h33f : errs =          31'b0000000000000000100000010000000; // D (0x00004080) 
10'h3f1 : errs =          31'b0000000000000000100000100000000; // D (0x00004100) 
10'h26d : errs =          31'b0000000000000000100001000000000; // D (0x00004200) 
10'h155 : errs =          31'b0000000000000000100010000000000; // D (0x00004400) 
10'h04c : errs =          31'b0000000000000000100100000000000; // D (0x00004800) 
10'h27e : errs =          31'b0000000000000000101000000000000; // D (0x00005000) 
10'h173 : errs =          31'b0000000000000000110000000000000; // D (0x00006000) 
10'h1a2 : errs =          31'b0000000000000000100000000000000; // S (0x00004000) 
//10'h2e6 : errs =          31'b0000000000000001100000000000000; // D (0x0000c000) 
//10'h043 : errs =          31'b0000000000000010100000000000000; // D (0x00014000) 
//10'h260 : errs =          31'b0000000000000100100000000000000; // D (0x00024000) 
//10'h14f : errs =          31'b0000000000001000100000000000000; // D (0x00044000) 
//10'h078 : errs =          31'b0000000000010000100000000000000; // D (0x00084000) 
//10'h216 : errs =          31'b0000000000100000100000000000000; // D (0x00104000) 
//10'h1a3 : errs =          31'b0000000001000000100000000000000; // D (0x00204000) 
//10'h1a0 : errs =          31'b0000000010000000100000000000000; // D (0x00404000) 
//10'h1a6 : errs =          31'b0000000100000000100000000000000; // D (0x00804000) 
//10'h1aa : errs =          31'b0000001000000000100000000000000; // D (0x01004000) 
//10'h1b2 : errs =          31'b0000010000000000100000000000000; // D (0x02004000) 
//10'h182 : errs =          31'b0000100000000000100000000000000; // D (0x04004000) 
//10'h1e2 : errs =          31'b0001000000000000100000000000000; // D (0x08004000) 
//10'h122 : errs =          31'b0010000000000000100000000000000; // D (0x10004000) 
//10'h0a2 : errs =          31'b0100000000000000100000000000000; // D (0x20004000) 
//10'h3a2 : errs =          31'b1000000000000000100000000000000; // D (0x40004000) 
10'h02d : errs =          31'b0000000000000001000000000000001; // D (0x00008001) 
10'h2ff : errs =          31'b0000000000000001000000000000010; // D (0x00008002) 
10'h032 : errs =          31'b0000000000000001000000000000100; // D (0x00008004) 
10'h2c1 : errs =          31'b0000000000000001000000000001000; // D (0x00008008) 
10'h04e : errs =          31'b0000000000000001000000000010000; // D (0x00008010) 
10'h239 : errs =          31'b0000000000000001000000000100000; // D (0x00008020) 
10'h1be : errs =          31'b0000000000000001000000001000000; // D (0x00008040) 
10'h1d9 : errs =          31'b0000000000000001000000010000000; // D (0x00008080) 
10'h117 : errs =          31'b0000000000000001000000100000000; // D (0x00008100) 
10'h08b : errs =          31'b0000000000000001000001000000000; // D (0x00008200) 
10'h3b3 : errs =          31'b0000000000000001000010000000000; // D (0x00008400) 
10'h2aa : errs =          31'b0000000000000001000100000000000; // D (0x00008800) 
10'h098 : errs =          31'b0000000000000001001000000000000; // D (0x00009000) 
10'h395 : errs =          31'b0000000000000001010000000000000; // D (0x0000a000) 
10'h2e6 : errs =          31'b0000000000000001100000000000000; // D (0x0000c000) 
10'h344 : errs =          31'b0000000000000001000000000000000; // S (0x00008000) 
//10'h2a5 : errs =          31'b0000000000000011000000000000000; // D (0x00018000) 
//10'h086 : errs =          31'b0000000000000101000000000000000; // D (0x00028000) 
//10'h3a9 : errs =          31'b0000000000001001000000000000000; // D (0x00048000) 
//10'h29e : errs =          31'b0000000000010001000000000000000; // D (0x00088000) 
//10'h0f0 : errs =          31'b0000000000100001000000000000000; // D (0x00108000) 
//10'h345 : errs =          31'b0000000001000001000000000000000; // D (0x00208000) 
//10'h346 : errs =          31'b0000000010000001000000000000000; // D (0x00408000) 
//10'h340 : errs =          31'b0000000100000001000000000000000; // D (0x00808000) 
//10'h34c : errs =          31'b0000001000000001000000000000000; // D (0x01008000) 
//10'h354 : errs =          31'b0000010000000001000000000000000; // D (0x02008000) 
//10'h364 : errs =          31'b0000100000000001000000000000000; // D (0x04008000) 
//10'h304 : errs =          31'b0001000000000001000000000000000; // D (0x08008000) 
//10'h3c4 : errs =          31'b0010000000000001000000000000000; // D (0x10008000) 
//10'h244 : errs =          31'b0100000000000001000000000000000; // D (0x20008000) 
//10'h144 : errs =          31'b1000000000000001000000000000000; // D (0x40008000) 
10'h288 : errs =          31'b0000000000000010000000000000001; // D (0x00010001) 
10'h05a : errs =          31'b0000000000000010000000000000010; // D (0x00010002) 
10'h297 : errs =          31'b0000000000000010000000000000100; // D (0x00010004) 
10'h064 : errs =          31'b0000000000000010000000000001000; // D (0x00010008) 
10'h2eb : errs =          31'b0000000000000010000000000010000; // D (0x00010010) 
10'h09c : errs =          31'b0000000000000010000000000100000; // D (0x00010020) 
10'h31b : errs =          31'b0000000000000010000000001000000; // D (0x00010040) 
10'h37c : errs =          31'b0000000000000010000000010000000; // D (0x00010080) 
10'h3b2 : errs =          31'b0000000000000010000000100000000; // D (0x00010100) 
10'h22e : errs =          31'b0000000000000010000001000000000; // D (0x00010200) 
10'h116 : errs =          31'b0000000000000010000010000000000; // D (0x00010400) 
10'h00f : errs =          31'b0000000000000010000100000000000; // D (0x00010800) 
10'h23d : errs =          31'b0000000000000010001000000000000; // D (0x00011000) 
10'h130 : errs =          31'b0000000000000010010000000000000; // D (0x00012000) 
10'h043 : errs =          31'b0000000000000010100000000000000; // D (0x00014000) 
10'h2a5 : errs =          31'b0000000000000011000000000000000; // D (0x00018000) 
10'h1e1 : errs =          31'b0000000000000010000000000000000; // S (0x00010000) 
//10'h223 : errs =          31'b0000000000000110000000000000000; // D (0x00030000) 
//10'h10c : errs =          31'b0000000000001010000000000000000; // D (0x00050000) 
//10'h03b : errs =          31'b0000000000010010000000000000000; // D (0x00090000) 
//10'h255 : errs =          31'b0000000000100010000000000000000; // D (0x00110000) 
//10'h1e0 : errs =          31'b0000000001000010000000000000000; // D (0x00210000) 
//10'h1e3 : errs =          31'b0000000010000010000000000000000; // D (0x00410000) 
//10'h1e5 : errs =          31'b0000000100000010000000000000000; // D (0x00810000) 
//10'h1e9 : errs =          31'b0000001000000010000000000000000; // D (0x01010000) 
//10'h1f1 : errs =          31'b0000010000000010000000000000000; // D (0x02010000) 
//10'h1c1 : errs =          31'b0000100000000010000000000000000; // D (0x04010000) 
//10'h1a1 : errs =          31'b0001000000000010000000000000000; // D (0x08010000) 
//10'h161 : errs =          31'b0010000000000010000000000000000; // D (0x10010000) 
//10'h0e1 : errs =          31'b0100000000000010000000000000000; // D (0x20010000) 
//10'h3e1 : errs =          31'b1000000000000010000000000000000; // D (0x40010000) 
10'h0ab : errs =          31'b0000000000000100000000000000001; // D (0x00020001) 
10'h279 : errs =          31'b0000000000000100000000000000010; // D (0x00020002) 
10'h0b4 : errs =          31'b0000000000000100000000000000100; // D (0x00020004) 
10'h247 : errs =          31'b0000000000000100000000000001000; // D (0x00020008) 
10'h0c8 : errs =          31'b0000000000000100000000000010000; // D (0x00020010) 
10'h2bf : errs =          31'b0000000000000100000000000100000; // D (0x00020020) 
10'h138 : errs =          31'b0000000000000100000000001000000; // D (0x00020040) 
10'h15f : errs =          31'b0000000000000100000000010000000; // D (0x00020080) 
10'h191 : errs =          31'b0000000000000100000000100000000; // D (0x00020100) 
10'h00d : errs =          31'b0000000000000100000001000000000; // D (0x00020200) 
10'h335 : errs =          31'b0000000000000100000010000000000; // D (0x00020400) 
10'h22c : errs =          31'b0000000000000100000100000000000; // D (0x00020800) 
10'h01e : errs =          31'b0000000000000100001000000000000; // D (0x00021000) 
10'h313 : errs =          31'b0000000000000100010000000000000; // D (0x00022000) 
10'h260 : errs =          31'b0000000000000100100000000000000; // D (0x00024000) 
10'h086 : errs =          31'b0000000000000101000000000000000; // D (0x00028000) 
10'h223 : errs =          31'b0000000000000110000000000000000; // D (0x00030000) 
10'h3c2 : errs =          31'b0000000000000100000000000000000; // S (0x00020000) 
//10'h32f : errs =          31'b0000000000001100000000000000000; // D (0x00060000) 
//10'h218 : errs =          31'b0000000000010100000000000000000; // D (0x000a0000) 
//10'h076 : errs =          31'b0000000000100100000000000000000; // D (0x00120000) 
//10'h3c3 : errs =          31'b0000000001000100000000000000000; // D (0x00220000) 
//10'h3c0 : errs =          31'b0000000010000100000000000000000; // D (0x00420000) 
//10'h3c6 : errs =          31'b0000000100000100000000000000000; // D (0x00820000) 
//10'h3ca : errs =          31'b0000001000000100000000000000000; // D (0x01020000) 
//10'h3d2 : errs =          31'b0000010000000100000000000000000; // D (0x02020000) 
//10'h3e2 : errs =          31'b0000100000000100000000000000000; // D (0x04020000) 
//10'h382 : errs =          31'b0001000000000100000000000000000; // D (0x08020000) 
//10'h342 : errs =          31'b0010000000000100000000000000000; // D (0x10020000) 
//10'h2c2 : errs =          31'b0100000000000100000000000000000; // D (0x20020000) 
//10'h1c2 : errs =          31'b1000000000000100000000000000000; // D (0x40020000) 
10'h384 : errs =          31'b0000000000001000000000000000001; // D (0x00040001) 
10'h156 : errs =          31'b0000000000001000000000000000010; // D (0x00040002) 
10'h39b : errs =          31'b0000000000001000000000000000100; // D (0x00040004) 
10'h168 : errs =          31'b0000000000001000000000000001000; // D (0x00040008) 
10'h3e7 : errs =          31'b0000000000001000000000000010000; // D (0x00040010) 
10'h190 : errs =          31'b0000000000001000000000000100000; // D (0x00040020) 
10'h217 : errs =          31'b0000000000001000000000001000000; // D (0x00040040) 
10'h270 : errs =          31'b0000000000001000000000010000000; // D (0x00040080) 
10'h2be : errs =          31'b0000000000001000000000100000000; // D (0x00040100) 
10'h322 : errs =          31'b0000000000001000000001000000000; // D (0x00040200) 
10'h01a : errs =          31'b0000000000001000000010000000000; // D (0x00040400) 
10'h103 : errs =          31'b0000000000001000000100000000000; // D (0x00040800) 
10'h331 : errs =          31'b0000000000001000001000000000000; // D (0x00041000) 
10'h03c : errs =          31'b0000000000001000010000000000000; // D (0x00042000) 
10'h14f : errs =          31'b0000000000001000100000000000000; // D (0x00044000) 
10'h3a9 : errs =          31'b0000000000001001000000000000000; // D (0x00048000) 
10'h10c : errs =          31'b0000000000001010000000000000000; // D (0x00050000) 
10'h32f : errs =          31'b0000000000001100000000000000000; // D (0x00060000) 
10'h0ed : errs =          31'b0000000000001000000000000000000; // S (0x00040000) 
//10'h137 : errs =          31'b0000000000011000000000000000000; // D (0x000c0000) 
//10'h359 : errs =          31'b0000000000101000000000000000000; // D (0x00140000) 
//10'h0ec : errs =          31'b0000000001001000000000000000000; // D (0x00240000) 
//10'h0ef : errs =          31'b0000000010001000000000000000000; // D (0x00440000) 
//10'h0e9 : errs =          31'b0000000100001000000000000000000; // D (0x00840000) 
//10'h0e5 : errs =          31'b0000001000001000000000000000000; // D (0x01040000) 
//10'h0fd : errs =          31'b0000010000001000000000000000000; // D (0x02040000) 
//10'h0cd : errs =          31'b0000100000001000000000000000000; // D (0x04040000) 
//10'h0ad : errs =          31'b0001000000001000000000000000000; // D (0x08040000) 
//10'h06d : errs =          31'b0010000000001000000000000000000; // D (0x10040000) 
//10'h1ed : errs =          31'b0100000000001000000000000000000; // D (0x20040000) 
//10'h2ed : errs =          31'b1000000000001000000000000000000; // D (0x40040000) 
10'h2b3 : errs =          31'b0000000000010000000000000000001; // D (0x00080001) 
10'h061 : errs =          31'b0000000000010000000000000000010; // D (0x00080002) 
10'h2ac : errs =          31'b0000000000010000000000000000100; // D (0x00080004) 
10'h05f : errs =          31'b0000000000010000000000000001000; // D (0x00080008) 
10'h2d0 : errs =          31'b0000000000010000000000000010000; // D (0x00080010) 
10'h0a7 : errs =          31'b0000000000010000000000000100000; // D (0x00080020) 
10'h320 : errs =          31'b0000000000010000000000001000000; // D (0x00080040) 
10'h347 : errs =          31'b0000000000010000000000010000000; // D (0x00080080) 
10'h389 : errs =          31'b0000000000010000000000100000000; // D (0x00080100) 
10'h215 : errs =          31'b0000000000010000000001000000000; // D (0x00080200) 
10'h12d : errs =          31'b0000000000010000000010000000000; // D (0x00080400) 
10'h034 : errs =          31'b0000000000010000000100000000000; // D (0x00080800) 
10'h206 : errs =          31'b0000000000010000001000000000000; // D (0x00081000) 
10'h10b : errs =          31'b0000000000010000010000000000000; // D (0x00082000) 
10'h078 : errs =          31'b0000000000010000100000000000000; // D (0x00084000) 
10'h29e : errs =          31'b0000000000010001000000000000000; // D (0x00088000) 
10'h03b : errs =          31'b0000000000010010000000000000000; // D (0x00090000) 
10'h218 : errs =          31'b0000000000010100000000000000000; // D (0x000a0000) 
10'h137 : errs =          31'b0000000000011000000000000000000; // D (0x000c0000) 
10'h1da : errs =          31'b0000000000010000000000000000000; // S (0x00080000) 
//10'h26e : errs =          31'b0000000000110000000000000000000; // D (0x00180000) 
//10'h1db : errs =          31'b0000000001010000000000000000000; // D (0x00280000) 
//10'h1d8 : errs =          31'b0000000010010000000000000000000; // D (0x00480000) 
//10'h1de : errs =          31'b0000000100010000000000000000000; // D (0x00880000) 
//10'h1d2 : errs =          31'b0000001000010000000000000000000; // D (0x01080000) 
//10'h1ca : errs =          31'b0000010000010000000000000000000; // D (0x02080000) 
//10'h1fa : errs =          31'b0000100000010000000000000000000; // D (0x04080000) 
//10'h19a : errs =          31'b0001000000010000000000000000000; // D (0x08080000) 
//10'h15a : errs =          31'b0010000000010000000000000000000; // D (0x10080000) 
//10'h0da : errs =          31'b0100000000010000000000000000000; // D (0x20080000) 
//10'h3da : errs =          31'b1000000000010000000000000000000; // D (0x40080000) 
10'h0dd : errs =          31'b0000000000100000000000000000001; // D (0x00100001) 
10'h20f : errs =          31'b0000000000100000000000000000010; // D (0x00100002) 
10'h0c2 : errs =          31'b0000000000100000000000000000100; // D (0x00100004) 
10'h231 : errs =          31'b0000000000100000000000000001000; // D (0x00100008) 
10'h0be : errs =          31'b0000000000100000000000000010000; // D (0x00100010) 
10'h2c9 : errs =          31'b0000000000100000000000000100000; // D (0x00100020) 
10'h14e : errs =          31'b0000000000100000000000001000000; // D (0x00100040) 
10'h129 : errs =          31'b0000000000100000000000010000000; // D (0x00100080) 
10'h1e7 : errs =          31'b0000000000100000000000100000000; // D (0x00100100) 
10'h07b : errs =          31'b0000000000100000000001000000000; // D (0x00100200) 
10'h343 : errs =          31'b0000000000100000000010000000000; // D (0x00100400) 
10'h25a : errs =          31'b0000000000100000000100000000000; // D (0x00100800) 
10'h068 : errs =          31'b0000000000100000001000000000000; // D (0x00101000) 
10'h365 : errs =          31'b0000000000100000010000000000000; // D (0x00102000) 
10'h216 : errs =          31'b0000000000100000100000000000000; // D (0x00104000) 
10'h0f0 : errs =          31'b0000000000100001000000000000000; // D (0x00108000) 
10'h255 : errs =          31'b0000000000100010000000000000000; // D (0x00110000) 
10'h076 : errs =          31'b0000000000100100000000000000000; // D (0x00120000) 
10'h359 : errs =          31'b0000000000101000000000000000000; // D (0x00140000) 
10'h26e : errs =          31'b0000000000110000000000000000000; // D (0x00180000) 
10'h3b4 : errs =          31'b0000000000100000000000000000000; // S (0x00100000) 
//10'h3b5 : errs =          31'b0000000001100000000000000000000; // D (0x00300000) 
//10'h3b6 : errs =          31'b0000000010100000000000000000000; // D (0x00500000) 
//10'h3b0 : errs =          31'b0000000100100000000000000000000; // D (0x00900000) 
//10'h3bc : errs =          31'b0000001000100000000000000000000; // D (0x01100000) 
//10'h3a4 : errs =          31'b0000010000100000000000000000000; // D (0x02100000) 
//10'h394 : errs =          31'b0000100000100000000000000000000; // D (0x04100000) 
//10'h3f4 : errs =          31'b0001000000100000000000000000000; // D (0x08100000) 
//10'h334 : errs =          31'b0010000000100000000000000000000; // D (0x10100000) 
//10'h2b4 : errs =          31'b0100000000100000000000000000000; // D (0x20100000) 
//10'h1b4 : errs =          31'b1000000000100000000000000000000; // D (0x40100000) 
10'h368 : errs =          31'b0000000001000000000000000000001; // D (0x00200001) 
10'h1ba : errs =          31'b0000000001000000000000000000010; // D (0x00200002) 
10'h377 : errs =          31'b0000000001000000000000000000100; // D (0x00200004) 
10'h184 : errs =          31'b0000000001000000000000000001000; // D (0x00200008) 
10'h30b : errs =          31'b0000000001000000000000000010000; // D (0x00200010) 
10'h17c : errs =          31'b0000000001000000000000000100000; // D (0x00200020) 
10'h2fb : errs =          31'b0000000001000000000000001000000; // D (0x00200040) 
10'h29c : errs =          31'b0000000001000000000000010000000; // D (0x00200080) 
10'h252 : errs =          31'b0000000001000000000000100000000; // D (0x00200100) 
10'h3ce : errs =          31'b0000000001000000000001000000000; // D (0x00200200) 
10'h0f6 : errs =          31'b0000000001000000000010000000000; // D (0x00200400) 
10'h1ef : errs =          31'b0000000001000000000100000000000; // D (0x00200800) 
10'h3dd : errs =          31'b0000000001000000001000000000000; // D (0x00201000) 
10'h0d0 : errs =          31'b0000000001000000010000000000000; // D (0x00202000) 
10'h1a3 : errs =          31'b0000000001000000100000000000000; // D (0x00204000) 
10'h345 : errs =          31'b0000000001000001000000000000000; // D (0x00208000) 
10'h1e0 : errs =          31'b0000000001000010000000000000000; // D (0x00210000) 
10'h3c3 : errs =          31'b0000000001000100000000000000000; // D (0x00220000) 
10'h0ec : errs =          31'b0000000001001000000000000000000; // D (0x00240000) 
10'h1db : errs =          31'b0000000001010000000000000000000; // D (0x00280000) 
10'h3b5 : errs =          31'b0000000001100000000000000000000; // D (0x00300000) 
10'h001 : errs =          31'b0000000001000000000000000000000; // S (0x00200000) 
//10'h003 : errs =          31'b0000000011000000000000000000000; // D (0x00600000) 
//10'h005 : errs =          31'b0000000101000000000000000000000; // D (0x00a00000) 
//10'h009 : errs =          31'b0000001001000000000000000000000; // D (0x01200000) 
//10'h011 : errs =          31'b0000010001000000000000000000000; // D (0x02200000) 
//10'h021 : errs =          31'b0000100001000000000000000000000; // D (0x04200000) 
//10'h041 : errs =          31'b0001000001000000000000000000000; // D (0x08200000) 
//10'h081 : errs =          31'b0010000001000000000000000000000; // D (0x10200000) 
//10'h101 : errs =          31'b0100000001000000000000000000000; // D (0x20200000) 
//10'h201 : errs =          31'b1000000001000000000000000000000; // D (0x40200000) 
10'h36b : errs =          31'b0000000010000000000000000000001; // D (0x00400001) 
10'h1b9 : errs =          31'b0000000010000000000000000000010; // D (0x00400002) 
10'h374 : errs =          31'b0000000010000000000000000000100; // D (0x00400004) 
10'h187 : errs =          31'b0000000010000000000000000001000; // D (0x00400008) 
10'h308 : errs =          31'b0000000010000000000000000010000; // D (0x00400010) 
10'h17f : errs =          31'b0000000010000000000000000100000; // D (0x00400020) 
10'h2f8 : errs =          31'b0000000010000000000000001000000; // D (0x00400040) 
10'h29f : errs =          31'b0000000010000000000000010000000; // D (0x00400080) 
10'h251 : errs =          31'b0000000010000000000000100000000; // D (0x00400100) 
10'h3cd : errs =          31'b0000000010000000000001000000000; // D (0x00400200) 
10'h0f5 : errs =          31'b0000000010000000000010000000000; // D (0x00400400) 
10'h1ec : errs =          31'b0000000010000000000100000000000; // D (0x00400800) 
10'h3de : errs =          31'b0000000010000000001000000000000; // D (0x00401000) 
10'h0d3 : errs =          31'b0000000010000000010000000000000; // D (0x00402000) 
10'h1a0 : errs =          31'b0000000010000000100000000000000; // D (0x00404000) 
10'h346 : errs =          31'b0000000010000001000000000000000; // D (0x00408000) 
10'h1e3 : errs =          31'b0000000010000010000000000000000; // D (0x00410000) 
10'h3c0 : errs =          31'b0000000010000100000000000000000; // D (0x00420000) 
10'h0ef : errs =          31'b0000000010001000000000000000000; // D (0x00440000) 
10'h1d8 : errs =          31'b0000000010010000000000000000000; // D (0x00480000) 
10'h3b6 : errs =          31'b0000000010100000000000000000000; // D (0x00500000) 
10'h003 : errs =          31'b0000000011000000000000000000000; // D (0x00600000) 
10'h002 : errs =          31'b0000000010000000000000000000000; // S (0x00400000) 
//10'h006 : errs =          31'b0000000110000000000000000000000; // D (0x00c00000) 
//10'h00a : errs =          31'b0000001010000000000000000000000; // D (0x01400000) 
//10'h012 : errs =          31'b0000010010000000000000000000000; // D (0x02400000) 
//10'h022 : errs =          31'b0000100010000000000000000000000; // D (0x04400000) 
//10'h042 : errs =          31'b0001000010000000000000000000000; // D (0x08400000) 
//10'h082 : errs =          31'b0010000010000000000000000000000; // D (0x10400000) 
//10'h102 : errs =          31'b0100000010000000000000000000000; // D (0x20400000) 
//10'h202 : errs =          31'b1000000010000000000000000000000; // D (0x40400000) 
10'h36d : errs =          31'b0000000100000000000000000000001; // D (0x00800001) 
10'h1bf : errs =          31'b0000000100000000000000000000010; // D (0x00800002) 
10'h372 : errs =          31'b0000000100000000000000000000100; // D (0x00800004) 
10'h181 : errs =          31'b0000000100000000000000000001000; // D (0x00800008) 
10'h30e : errs =          31'b0000000100000000000000000010000; // D (0x00800010) 
10'h179 : errs =          31'b0000000100000000000000000100000; // D (0x00800020) 
10'h2fe : errs =          31'b0000000100000000000000001000000; // D (0x00800040) 
10'h299 : errs =          31'b0000000100000000000000010000000; // D (0x00800080) 
10'h257 : errs =          31'b0000000100000000000000100000000; // D (0x00800100) 
10'h3cb : errs =          31'b0000000100000000000001000000000; // D (0x00800200) 
10'h0f3 : errs =          31'b0000000100000000000010000000000; // D (0x00800400) 
10'h1ea : errs =          31'b0000000100000000000100000000000; // D (0x00800800) 
10'h3d8 : errs =          31'b0000000100000000001000000000000; // D (0x00801000) 
10'h0d5 : errs =          31'b0000000100000000010000000000000; // D (0x00802000) 
10'h1a6 : errs =          31'b0000000100000000100000000000000; // D (0x00804000) 
10'h340 : errs =          31'b0000000100000001000000000000000; // D (0x00808000) 
10'h1e5 : errs =          31'b0000000100000010000000000000000; // D (0x00810000) 
10'h3c6 : errs =          31'b0000000100000100000000000000000; // D (0x00820000) 
10'h0e9 : errs =          31'b0000000100001000000000000000000; // D (0x00840000) 
10'h1de : errs =          31'b0000000100010000000000000000000; // D (0x00880000) 
10'h3b0 : errs =          31'b0000000100100000000000000000000; // D (0x00900000) 
10'h005 : errs =          31'b0000000101000000000000000000000; // D (0x00a00000) 
10'h006 : errs =          31'b0000000110000000000000000000000; // D (0x00c00000) 
10'h004 : errs =          31'b0000000100000000000000000000000; // S (0x00800000) 
//10'h00c : errs =          31'b0000001100000000000000000000000; // D (0x01800000) 
//10'h014 : errs =          31'b0000010100000000000000000000000; // D (0x02800000) 
//10'h024 : errs =          31'b0000100100000000000000000000000; // D (0x04800000) 
//10'h044 : errs =          31'b0001000100000000000000000000000; // D (0x08800000) 
//10'h084 : errs =          31'b0010000100000000000000000000000; // D (0x10800000) 
//10'h104 : errs =          31'b0100000100000000000000000000000; // D (0x20800000) 
//10'h204 : errs =          31'b1000000100000000000000000000000; // D (0x40800000) 
10'h361 : errs =          31'b0000001000000000000000000000001; // D (0x01000001) 
10'h1b3 : errs =          31'b0000001000000000000000000000010; // D (0x01000002) 
10'h37e : errs =          31'b0000001000000000000000000000100; // D (0x01000004) 
10'h18d : errs =          31'b0000001000000000000000000001000; // D (0x01000008) 
10'h302 : errs =          31'b0000001000000000000000000010000; // D (0x01000010) 
10'h175 : errs =          31'b0000001000000000000000000100000; // D (0x01000020) 
10'h2f2 : errs =          31'b0000001000000000000000001000000; // D (0x01000040) 
10'h295 : errs =          31'b0000001000000000000000010000000; // D (0x01000080) 
10'h25b : errs =          31'b0000001000000000000000100000000; // D (0x01000100) 
10'h3c7 : errs =          31'b0000001000000000000001000000000; // D (0x01000200) 
10'h0ff : errs =          31'b0000001000000000000010000000000; // D (0x01000400) 
10'h1e6 : errs =          31'b0000001000000000000100000000000; // D (0x01000800) 
10'h3d4 : errs =          31'b0000001000000000001000000000000; // D (0x01001000) 
10'h0d9 : errs =          31'b0000001000000000010000000000000; // D (0x01002000) 
10'h1aa : errs =          31'b0000001000000000100000000000000; // D (0x01004000) 
10'h34c : errs =          31'b0000001000000001000000000000000; // D (0x01008000) 
10'h1e9 : errs =          31'b0000001000000010000000000000000; // D (0x01010000) 
10'h3ca : errs =          31'b0000001000000100000000000000000; // D (0x01020000) 
10'h0e5 : errs =          31'b0000001000001000000000000000000; // D (0x01040000) 
10'h1d2 : errs =          31'b0000001000010000000000000000000; // D (0x01080000) 
10'h3bc : errs =          31'b0000001000100000000000000000000; // D (0x01100000) 
10'h009 : errs =          31'b0000001001000000000000000000000; // D (0x01200000) 
10'h00a : errs =          31'b0000001010000000000000000000000; // D (0x01400000) 
10'h00c : errs =          31'b0000001100000000000000000000000; // D (0x01800000) 
10'h008 : errs =          31'b0000001000000000000000000000000; // S (0x01000000) 
//10'h018 : errs =          31'b0000011000000000000000000000000; // D (0x03000000) 
//10'h028 : errs =          31'b0000101000000000000000000000000; // D (0x05000000) 
//10'h048 : errs =          31'b0001001000000000000000000000000; // D (0x09000000) 
//10'h088 : errs =          31'b0010001000000000000000000000000; // D (0x11000000) 
//10'h108 : errs =          31'b0100001000000000000000000000000; // D (0x21000000) 
//10'h208 : errs =          31'b1000001000000000000000000000000; // D (0x41000000) 
10'h379 : errs =          31'b0000010000000000000000000000001; // D (0x02000001) 
10'h1ab : errs =          31'b0000010000000000000000000000010; // D (0x02000002) 
10'h366 : errs =          31'b0000010000000000000000000000100; // D (0x02000004) 
10'h195 : errs =          31'b0000010000000000000000000001000; // D (0x02000008) 
10'h31a : errs =          31'b0000010000000000000000000010000; // D (0x02000010) 
10'h16d : errs =          31'b0000010000000000000000000100000; // D (0x02000020) 
10'h2ea : errs =          31'b0000010000000000000000001000000; // D (0x02000040) 
10'h28d : errs =          31'b0000010000000000000000010000000; // D (0x02000080) 
10'h243 : errs =          31'b0000010000000000000000100000000; // D (0x02000100) 
10'h3df : errs =          31'b0000010000000000000001000000000; // D (0x02000200) 
10'h0e7 : errs =          31'b0000010000000000000010000000000; // D (0x02000400) 
10'h1fe : errs =          31'b0000010000000000000100000000000; // D (0x02000800) 
10'h3cc : errs =          31'b0000010000000000001000000000000; // D (0x02001000) 
10'h0c1 : errs =          31'b0000010000000000010000000000000; // D (0x02002000) 
10'h1b2 : errs =          31'b0000010000000000100000000000000; // D (0x02004000) 
10'h354 : errs =          31'b0000010000000001000000000000000; // D (0x02008000) 
10'h1f1 : errs =          31'b0000010000000010000000000000000; // D (0x02010000) 
10'h3d2 : errs =          31'b0000010000000100000000000000000; // D (0x02020000) 
10'h0fd : errs =          31'b0000010000001000000000000000000; // D (0x02040000) 
10'h1ca : errs =          31'b0000010000010000000000000000000; // D (0x02080000) 
10'h3a4 : errs =          31'b0000010000100000000000000000000; // D (0x02100000) 
10'h011 : errs =          31'b0000010001000000000000000000000; // D (0x02200000) 
10'h012 : errs =          31'b0000010010000000000000000000000; // D (0x02400000) 
10'h014 : errs =          31'b0000010100000000000000000000000; // D (0x02800000) 
10'h018 : errs =          31'b0000011000000000000000000000000; // D (0x03000000) 
10'h010 : errs =          31'b0000010000000000000000000000000; // S (0x02000000) 
//10'h030 : errs =          31'b0000110000000000000000000000000; // D (0x06000000) 
//10'h050 : errs =          31'b0001010000000000000000000000000; // D (0x0a000000) 
//10'h090 : errs =          31'b0010010000000000000000000000000; // D (0x12000000) 
//10'h110 : errs =          31'b0100010000000000000000000000000; // D (0x22000000) 
//10'h210 : errs =          31'b1000010000000000000000000000000; // D (0x42000000) 
10'h349 : errs =          31'b0000100000000000000000000000001; // D (0x04000001) 
10'h19b : errs =          31'b0000100000000000000000000000010; // D (0x04000002) 
10'h356 : errs =          31'b0000100000000000000000000000100; // D (0x04000004) 
10'h1a5 : errs =          31'b0000100000000000000000000001000; // D (0x04000008) 
10'h32a : errs =          31'b0000100000000000000000000010000; // D (0x04000010) 
10'h15d : errs =          31'b0000100000000000000000000100000; // D (0x04000020) 
10'h2da : errs =          31'b0000100000000000000000001000000; // D (0x04000040) 
10'h2bd : errs =          31'b0000100000000000000000010000000; // D (0x04000080) 
10'h273 : errs =          31'b0000100000000000000000100000000; // D (0x04000100) 
10'h3ef : errs =          31'b0000100000000000000001000000000; // D (0x04000200) 
10'h0d7 : errs =          31'b0000100000000000000010000000000; // D (0x04000400) 
10'h1ce : errs =          31'b0000100000000000000100000000000; // D (0x04000800) 
10'h3fc : errs =          31'b0000100000000000001000000000000; // D (0x04001000) 
10'h0f1 : errs =          31'b0000100000000000010000000000000; // D (0x04002000) 
10'h182 : errs =          31'b0000100000000000100000000000000; // D (0x04004000) 
10'h364 : errs =          31'b0000100000000001000000000000000; // D (0x04008000) 
10'h1c1 : errs =          31'b0000100000000010000000000000000; // D (0x04010000) 
10'h3e2 : errs =          31'b0000100000000100000000000000000; // D (0x04020000) 
10'h0cd : errs =          31'b0000100000001000000000000000000; // D (0x04040000) 
10'h1fa : errs =          31'b0000100000010000000000000000000; // D (0x04080000) 
10'h394 : errs =          31'b0000100000100000000000000000000; // D (0x04100000) 
10'h021 : errs =          31'b0000100001000000000000000000000; // D (0x04200000) 
10'h022 : errs =          31'b0000100010000000000000000000000; // D (0x04400000) 
10'h024 : errs =          31'b0000100100000000000000000000000; // D (0x04800000) 
10'h028 : errs =          31'b0000101000000000000000000000000; // D (0x05000000) 
10'h030 : errs =          31'b0000110000000000000000000000000; // D (0x06000000) 
10'h020 : errs =          31'b0000100000000000000000000000000; // S (0x04000000) 
//10'h060 : errs =          31'b0001100000000000000000000000000; // D (0x0c000000) 
//10'h0a0 : errs =          31'b0010100000000000000000000000000; // D (0x14000000) 
//10'h120 : errs =          31'b0100100000000000000000000000000; // D (0x24000000) 
//10'h220 : errs =          31'b1000100000000000000000000000000; // D (0x44000000) 
10'h329 : errs =          31'b0001000000000000000000000000001; // D (0x08000001) 
10'h1fb : errs =          31'b0001000000000000000000000000010; // D (0x08000002) 
10'h336 : errs =          31'b0001000000000000000000000000100; // D (0x08000004) 
10'h1c5 : errs =          31'b0001000000000000000000000001000; // D (0x08000008) 
10'h34a : errs =          31'b0001000000000000000000000010000; // D (0x08000010) 
10'h13d : errs =          31'b0001000000000000000000000100000; // D (0x08000020) 
10'h2ba : errs =          31'b0001000000000000000000001000000; // D (0x08000040) 
10'h2dd : errs =          31'b0001000000000000000000010000000; // D (0x08000080) 
10'h213 : errs =          31'b0001000000000000000000100000000; // D (0x08000100) 
10'h38f : errs =          31'b0001000000000000000001000000000; // D (0x08000200) 
10'h0b7 : errs =          31'b0001000000000000000010000000000; // D (0x08000400) 
10'h1ae : errs =          31'b0001000000000000000100000000000; // D (0x08000800) 
10'h39c : errs =          31'b0001000000000000001000000000000; // D (0x08001000) 
10'h091 : errs =          31'b0001000000000000010000000000000; // D (0x08002000) 
10'h1e2 : errs =          31'b0001000000000000100000000000000; // D (0x08004000) 
10'h304 : errs =          31'b0001000000000001000000000000000; // D (0x08008000) 
10'h1a1 : errs =          31'b0001000000000010000000000000000; // D (0x08010000) 
10'h382 : errs =          31'b0001000000000100000000000000000; // D (0x08020000) 
10'h0ad : errs =          31'b0001000000001000000000000000000; // D (0x08040000) 
10'h19a : errs =          31'b0001000000010000000000000000000; // D (0x08080000) 
10'h3f4 : errs =          31'b0001000000100000000000000000000; // D (0x08100000) 
10'h041 : errs =          31'b0001000001000000000000000000000; // D (0x08200000) 
10'h042 : errs =          31'b0001000010000000000000000000000; // D (0x08400000) 
10'h044 : errs =          31'b0001000100000000000000000000000; // D (0x08800000) 
10'h048 : errs =          31'b0001001000000000000000000000000; // D (0x09000000) 
10'h050 : errs =          31'b0001010000000000000000000000000; // D (0x0a000000) 
10'h060 : errs =          31'b0001100000000000000000000000000; // D (0x0c000000) 
10'h040 : errs =          31'b0001000000000000000000000000000; // S (0x08000000) 
//10'h0c0 : errs =          31'b0011000000000000000000000000000; // D (0x18000000) 
//10'h140 : errs =          31'b0101000000000000000000000000000; // D (0x28000000) 
//10'h240 : errs =          31'b1001000000000000000000000000000; // D (0x48000000) 
10'h3e9 : errs =          31'b0010000000000000000000000000001; // D (0x10000001) 
10'h13b : errs =          31'b0010000000000000000000000000010; // D (0x10000002) 
10'h3f6 : errs =          31'b0010000000000000000000000000100; // D (0x10000004) 
10'h105 : errs =          31'b0010000000000000000000000001000; // D (0x10000008) 
10'h38a : errs =          31'b0010000000000000000000000010000; // D (0x10000010) 
10'h1fd : errs =          31'b0010000000000000000000000100000; // D (0x10000020) 
10'h27a : errs =          31'b0010000000000000000000001000000; // D (0x10000040) 
10'h21d : errs =          31'b0010000000000000000000010000000; // D (0x10000080) 
10'h2d3 : errs =          31'b0010000000000000000000100000000; // D (0x10000100) 
10'h34f : errs =          31'b0010000000000000000001000000000; // D (0x10000200) 
10'h077 : errs =          31'b0010000000000000000010000000000; // D (0x10000400) 
10'h16e : errs =          31'b0010000000000000000100000000000; // D (0x10000800) 
10'h35c : errs =          31'b0010000000000000001000000000000; // D (0x10001000) 
10'h051 : errs =          31'b0010000000000000010000000000000; // D (0x10002000) 
10'h122 : errs =          31'b0010000000000000100000000000000; // D (0x10004000) 
10'h3c4 : errs =          31'b0010000000000001000000000000000; // D (0x10008000) 
10'h161 : errs =          31'b0010000000000010000000000000000; // D (0x10010000) 
10'h342 : errs =          31'b0010000000000100000000000000000; // D (0x10020000) 
10'h06d : errs =          31'b0010000000001000000000000000000; // D (0x10040000) 
10'h15a : errs =          31'b0010000000010000000000000000000; // D (0x10080000) 
10'h334 : errs =          31'b0010000000100000000000000000000; // D (0x10100000) 
10'h081 : errs =          31'b0010000001000000000000000000000; // D (0x10200000) 
10'h082 : errs =          31'b0010000010000000000000000000000; // D (0x10400000) 
10'h084 : errs =          31'b0010000100000000000000000000000; // D (0x10800000) 
10'h088 : errs =          31'b0010001000000000000000000000000; // D (0x11000000) 
10'h090 : errs =          31'b0010010000000000000000000000000; // D (0x12000000) 
10'h0a0 : errs =          31'b0010100000000000000000000000000; // D (0x14000000) 
10'h0c0 : errs =          31'b0011000000000000000000000000000; // D (0x18000000) 
10'h080 : errs =          31'b0010000000000000000000000000000; // S (0x10000000) 
//10'h180 : errs =          31'b0110000000000000000000000000000; // D (0x30000000) 
//10'h280 : errs =          31'b1010000000000000000000000000000; // D (0x50000000) 
10'h269 : errs =          31'b0100000000000000000000000000001; // D (0x20000001) 
10'h0bb : errs =          31'b0100000000000000000000000000010; // D (0x20000002) 
10'h276 : errs =          31'b0100000000000000000000000000100; // D (0x20000004) 
10'h085 : errs =          31'b0100000000000000000000000001000; // D (0x20000008) 
10'h20a : errs =          31'b0100000000000000000000000010000; // D (0x20000010) 
10'h07d : errs =          31'b0100000000000000000000000100000; // D (0x20000020) 
10'h3fa : errs =          31'b0100000000000000000000001000000; // D (0x20000040) 
10'h39d : errs =          31'b0100000000000000000000010000000; // D (0x20000080) 
10'h353 : errs =          31'b0100000000000000000000100000000; // D (0x20000100) 
10'h2cf : errs =          31'b0100000000000000000001000000000; // D (0x20000200) 
10'h1f7 : errs =          31'b0100000000000000000010000000000; // D (0x20000400) 
10'h0ee : errs =          31'b0100000000000000000100000000000; // D (0x20000800) 
10'h2dc : errs =          31'b0100000000000000001000000000000; // D (0x20001000) 
10'h1d1 : errs =          31'b0100000000000000010000000000000; // D (0x20002000) 
10'h0a2 : errs =          31'b0100000000000000100000000000000; // D (0x20004000) 
10'h244 : errs =          31'b0100000000000001000000000000000; // D (0x20008000) 
10'h0e1 : errs =          31'b0100000000000010000000000000000; // D (0x20010000) 
10'h2c2 : errs =          31'b0100000000000100000000000000000; // D (0x20020000) 
10'h1ed : errs =          31'b0100000000001000000000000000000; // D (0x20040000) 
10'h0da : errs =          31'b0100000000010000000000000000000; // D (0x20080000) 
10'h2b4 : errs =          31'b0100000000100000000000000000000; // D (0x20100000) 
10'h101 : errs =          31'b0100000001000000000000000000000; // D (0x20200000) 
10'h102 : errs =          31'b0100000010000000000000000000000; // D (0x20400000) 
10'h104 : errs =          31'b0100000100000000000000000000000; // D (0x20800000) 
10'h108 : errs =          31'b0100001000000000000000000000000; // D (0x21000000) 
10'h110 : errs =          31'b0100010000000000000000000000000; // D (0x22000000) 
10'h120 : errs =          31'b0100100000000000000000000000000; // D (0x24000000) 
10'h140 : errs =          31'b0101000000000000000000000000000; // D (0x28000000) 
10'h180 : errs =          31'b0110000000000000000000000000000; // D (0x30000000) 
10'h100 : errs =          31'b0100000000000000000000000000000; // S (0x20000000) 
//10'h300 : errs =          31'b1100000000000000000000000000000; // D (0x60000000) 
10'h169 : errs =          31'b1000000000000000000000000000001; // D (0x40000001) 
10'h3bb : errs =          31'b1000000000000000000000000000010; // D (0x40000002) 
10'h176 : errs =          31'b1000000000000000000000000000100; // D (0x40000004) 
10'h385 : errs =          31'b1000000000000000000000000001000; // D (0x40000008) 
10'h10a : errs =          31'b1000000000000000000000000010000; // D (0x40000010) 
10'h37d : errs =          31'b1000000000000000000000000100000; // D (0x40000020) 
10'h0fa : errs =          31'b1000000000000000000000001000000; // D (0x40000040) 
10'h09d : errs =          31'b1000000000000000000000010000000; // D (0x40000080) 
10'h053 : errs =          31'b1000000000000000000000100000000; // D (0x40000100) 
10'h1cf : errs =          31'b1000000000000000000001000000000; // D (0x40000200) 
10'h2f7 : errs =          31'b1000000000000000000010000000000; // D (0x40000400) 
10'h3ee : errs =          31'b1000000000000000000100000000000; // D (0x40000800) 
10'h1dc : errs =          31'b1000000000000000001000000000000; // D (0x40001000) 
10'h2d1 : errs =          31'b1000000000000000010000000000000; // D (0x40002000) 
10'h3a2 : errs =          31'b1000000000000000100000000000000; // D (0x40004000) 
10'h144 : errs =          31'b1000000000000001000000000000000; // D (0x40008000) 
10'h3e1 : errs =          31'b1000000000000010000000000000000; // D (0x40010000) 
10'h1c2 : errs =          31'b1000000000000100000000000000000; // D (0x40020000) 
10'h2ed : errs =          31'b1000000000001000000000000000000; // D (0x40040000) 
10'h3da : errs =          31'b1000000000010000000000000000000; // D (0x40080000) 
10'h1b4 : errs =          31'b1000000000100000000000000000000; // D (0x40100000) 
10'h201 : errs =          31'b1000000001000000000000000000000; // D (0x40200000) 
10'h202 : errs =          31'b1000000010000000000000000000000; // D (0x40400000) 
10'h204 : errs =          31'b1000000100000000000000000000000; // D (0x40800000) 
10'h208 : errs =          31'b1000001000000000000000000000000; // D (0x41000000) 
10'h210 : errs =          31'b1000010000000000000000000000000; // D (0x42000000) 
10'h220 : errs =          31'b1000100000000000000000000000000; // D (0x44000000) 
10'h240 : errs =          31'b1001000000000000000000000000000; // D (0x48000000) 
10'h280 : errs =          31'b1010000000000000000000000000000; // D (0x50000000) 
10'h300 : errs =          31'b1100000000000000000000000000000; // D (0x60000000) 
10'h200 : errs =          31'b1000000000000000000000000000000; // S (0x40000000) 	 
default : errs = {(31){1'b0}};     
 endcase	

// Num of errs. =         961. Single =          31. Double =         930

 fn_err_pat_dcd_gf5_rom = errs; 
 
end						
endfunction // fn_err_pat_dcd_gf5_rom				
